module LERP(
  input  [16:0] io_samples_0,
  input  [16:0] io_samples_1,
  input  [9:0]  io_index,
  output [16:0] io_out
);

  wire [17:0] slope =
    18'({io_samples_1[16], io_samples_1} - {io_samples_0[16], io_samples_0});
  wire [25:0] _offset_T_1 = 26'({{8{slope[17]}}, slope} * {16'h0, io_index});
  assign io_out = 17'(_offset_T_1[25:9] + io_samples_0);
endmodule

