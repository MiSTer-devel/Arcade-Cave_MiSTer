module ReadCache_3(
  input         clock,
  input         reset,
  input         io_enable,
  input         io_in_rd,
  input  [31:0] io_in_addr,
  output [63:0] io_in_dout,
  output        io_in_wait_n,
  output        io_in_valid,
  output        io_out_rd,
  output [24:0] io_out_addr,
  input  [15:0] io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid
);

  wire [15:0] nextCacheEntry_line_words_3;
  wire [15:0] nextCacheEntry_line_words_2;
  wire [15:0] nextCacheEntry_line_words_1;
  wire [15:0] nextCacheEntry_line_words_0;
  wire [26:0] nextCacheEntry_tag;
  wire        nextCacheEntry_dirty;
  wire        nextCacheEntry_valid;
  wire [2:0]  _cacheEntryMemB_ext_R0_addr;
  wire        _cacheEntryMemB_ext_R0_en = 1'h1;
  wire        _cacheEntryMemB_ext_W0_en;
  wire [92:0] _cacheEntryMemB_ext_R0_data;
  wire [2:0]  _cacheEntryMemA_ext_R0_addr;
  wire        _cacheEntryMemA_ext_R0_en = 1'h1;
  wire        _cacheEntryMemA_ext_W0_en;
  wire [92:0] _cacheEntryMemA_ext_R0_data;
  reg  [2:0]  stateReg;
  reg         requestReg_rd;
  reg  [26:0] requestReg_addr_tag;
  reg  [2:0]  requestReg_addr_index;
  reg  [1:0]  requestReg_addr_offset;
  reg  [63:0] doutReg;
  reg         validReg;
  reg  [7:0]  lruReg;
  reg         wayReg;
  wire [92:0] _GEN =
    {nextCacheEntry_valid,
     nextCacheEntry_dirty,
     nextCacheEntry_tag,
     nextCacheEntry_line_words_3,
     nextCacheEntry_line_words_2,
     nextCacheEntry_line_words_1,
     nextCacheEntry_line_words_0};
  wire        _io_debug_check_T = stateReg == 3'h2;
  reg         cacheEntryReg_valid;
  reg         cacheEntryReg_dirty;
  reg  [26:0] cacheEntryReg_tag;
  reg  [15:0] cacheEntryReg_line_words_0;
  reg  [15:0] cacheEntryReg_line_words_1;
  reg  [15:0] cacheEntryReg_line_words_2;
  reg  [15:0] cacheEntryReg_line_words_3;
  wire        _io_debug_write_T = stateReg == 3'h5;
  assign nextCacheEntry_valid = _io_debug_write_T & cacheEntryReg_valid;
  assign nextCacheEntry_dirty = _io_debug_write_T & cacheEntryReg_dirty;
  assign nextCacheEntry_tag = _io_debug_write_T ? cacheEntryReg_tag : 27'h0;
  assign nextCacheEntry_line_words_0 =
    _io_debug_write_T ? cacheEntryReg_line_words_0 : 16'h0;
  assign nextCacheEntry_line_words_1 =
    _io_debug_write_T ? cacheEntryReg_line_words_1 : 16'h0;
  assign nextCacheEntry_line_words_2 =
    _io_debug_write_T ? cacheEntryReg_line_words_2 : 16'h0;
  assign nextCacheEntry_line_words_3 =
    _io_debug_write_T ? cacheEntryReg_line_words_3 : 16'h0;
  wire        _GEN_0 = stateReg == 3'h0;
  wire        _io_debug_fillWait_T = stateReg == 3'h4;
  wire        burstCounterEnable = _io_debug_fillWait_T & io_out_valid;
  reg  [2:0]  initCounter;
  reg  [1:0]  burstCounter;
  wire        _io_debug_idle_T = stateReg == 3'h1;
  wire        start = io_enable & io_in_rd & _io_debug_idle_T;
  wire        hitA =
    _cacheEntryMemA_ext_R0_data[92]
    & _cacheEntryMemA_ext_R0_data[90:64] == requestReg_addr_tag;
  wire        hit =
    hitA | _cacheEntryMemB_ext_R0_data[92]
    & _cacheEntryMemB_ext_R0_data[90:64] == requestReg_addr_tag;
  wire [7:0]  _nextWay_T = lruReg >> io_in_addr[5:3];
  wire        _nextWay_T_2 = start ? _nextWay_T[0] : wayReg;
  wire        _GEN_1 = _io_debug_check_T & hit;
  wire        _GEN_2 = _GEN_0 | _io_debug_idle_T;
  wire        _GEN_3 = _GEN_2 | ~_GEN_1;
  wire        nextWay = _GEN_3 ? _nextWay_T_2 : ~hitA;
  reg  [2:0]  casez_tmp;
  always @(*) begin
    casez (stateReg)
      3'b000:
        casez_tmp = _GEN_0 & (&initCounter) ? 3'h1 : stateReg;
      3'b001:
        casez_tmp = start ? 3'h2 : stateReg;
      3'b010:
        casez_tmp = {1'h0, ~hit, 1'h1};
      3'b011:
        casez_tmp = io_out_wait_n ? 3'h4 : stateReg;
      3'b100:
        casez_tmp = burstCounterEnable & (&burstCounter) ? 3'h5 : stateReg;
      3'b101:
        casez_tmp = 3'h1;
      3'b110:
        casez_tmp = stateReg;
      default:
        casez_tmp = stateReg;
    endcase
  end // always @(*)
  wire [7:0]  _GEN_4 = {5'h0, requestReg_addr_index};
  wire [7:0]  _lruReg_T = 8'h1 << _GEN_4;
  wire [7:0]  _lruReg_T_7 = 8'h1 << _GEN_4;
  wire [7:0]  _lruReg_T_12 = wayReg ? ~(~lruReg | _lruReg_T_7) : lruReg | _lruReg_T_7;
  wire [7:0]  _lruReg_T_5 = hitA ? lruReg | _lruReg_T : ~(~lruReg | _lruReg_T);
  wire        _GEN_5 = _io_debug_fillWait_T & io_out_valid;
  wire [1:0]  _n_T = 2'(requestReg_addr_offset + burstCounter);
  wire        _GEN_6 = _n_T == 2'h0;
  wire        _GEN_7 = _n_T == 2'h1;
  wire        _GEN_8 = _n_T == 2'h2;
  wire [15:0] entry_line_words_0 = _GEN_6 ? io_out_dout : cacheEntryReg_line_words_0;
  wire [15:0] entry_line_words_1 = _GEN_7 ? io_out_dout : cacheEntryReg_line_words_1;
  wire [15:0] entry_line_words_2 = _GEN_8 ? io_out_dout : cacheEntryReg_line_words_2;
  wire [15:0] entry_line_words_3 = (&_n_T) ? io_out_dout : cacheEntryReg_line_words_3;
  wire        _cacheEntryReg_T_valid =
    nextWay ? _cacheEntryMemB_ext_R0_data[92] : _cacheEntryMemA_ext_R0_data[92];
  wire        _GEN_9 = _io_debug_check_T ? _cacheEntryReg_T_valid : cacheEntryReg_valid;
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 3'h0;
      initCounter <= 3'h0;
      burstCounter <= 2'h0;
    end
    else begin
      stateReg <= casez_tmp;
      if (_GEN_0)
        initCounter <= 3'(initCounter + 3'h1);
      if (burstCounterEnable)
        burstCounter <= 2'(burstCounter + 2'h1);
    end
    if (start) begin
      requestReg_rd <= io_in_rd;
      requestReg_addr_tag <= {1'h0, io_in_addr[31:6]};
      requestReg_addr_index <= io_in_addr[5:3];
      requestReg_addr_offset <= io_in_addr[2:1];
    end
    if (_GEN_3) begin
      if (_GEN_5)
        doutReg <=
          {entry_line_words_0[7:0],
           entry_line_words_0[15:8],
           entry_line_words_1[7:0],
           entry_line_words_1[15:8],
           entry_line_words_2[7:0],
           entry_line_words_2[15:8],
           entry_line_words_3[7:0],
           entry_line_words_3[15:8]};
    end
    else
      doutReg <=
        hitA
          ? {_cacheEntryMemA_ext_R0_data[7:0],
             _cacheEntryMemA_ext_R0_data[15:8],
             _cacheEntryMemA_ext_R0_data[23:16],
             _cacheEntryMemA_ext_R0_data[31:24],
             _cacheEntryMemA_ext_R0_data[39:32],
             _cacheEntryMemA_ext_R0_data[47:40],
             _cacheEntryMemA_ext_R0_data[55:48],
             _cacheEntryMemA_ext_R0_data[63:56]}
          : {_cacheEntryMemB_ext_R0_data[7:0],
             _cacheEntryMemB_ext_R0_data[15:8],
             _cacheEntryMemB_ext_R0_data[23:16],
             _cacheEntryMemB_ext_R0_data[31:24],
             _cacheEntryMemB_ext_R0_data[39:32],
             _cacheEntryMemB_ext_R0_data[47:40],
             _cacheEntryMemB_ext_R0_data[55:48],
             _cacheEntryMemB_ext_R0_data[63:56]};
    validReg <= ~_GEN_2 & _GEN_1 | _GEN_5 & requestReg_rd & (&burstCounter);
    if (_GEN_2 | ~_io_debug_check_T) begin
    end
    else
      lruReg <= hit ? _lruReg_T_5 : _lruReg_T_12;
    if (_GEN_3) begin
      if (start)
        wayReg <= _nextWay_T[0];
    end
    else
      wayReg <= ~hitA;
    cacheEntryReg_valid <= _GEN_5 | _GEN_9;
    if (_GEN_5 | ~_io_debug_check_T) begin
    end
    else
      cacheEntryReg_dirty <=
        nextWay ? _cacheEntryMemB_ext_R0_data[91] : _cacheEntryMemA_ext_R0_data[91];
    if (_GEN_5) begin
      cacheEntryReg_tag <= requestReg_addr_tag;
      if (_GEN_6)
        cacheEntryReg_line_words_0 <= io_out_dout;
      if (_GEN_7)
        cacheEntryReg_line_words_1 <= io_out_dout;
      if (_GEN_8)
        cacheEntryReg_line_words_2 <= io_out_dout;
      if (&_n_T)
        cacheEntryReg_line_words_3 <= io_out_dout;
    end
    else if (_io_debug_check_T) begin
      cacheEntryReg_tag <=
        nextWay ? _cacheEntryMemB_ext_R0_data[90:64] : _cacheEntryMemA_ext_R0_data[90:64];
      cacheEntryReg_line_words_0 <=
        nextWay ? _cacheEntryMemB_ext_R0_data[15:0] : _cacheEntryMemA_ext_R0_data[15:0];
      cacheEntryReg_line_words_1 <=
        nextWay ? _cacheEntryMemB_ext_R0_data[31:16] : _cacheEntryMemA_ext_R0_data[31:16];
      cacheEntryReg_line_words_2 <=
        nextWay ? _cacheEntryMemB_ext_R0_data[47:32] : _cacheEntryMemA_ext_R0_data[47:32];
      cacheEntryReg_line_words_3 <=
        nextWay ? _cacheEntryMemB_ext_R0_data[63:48] : _cacheEntryMemA_ext_R0_data[63:48];
    end
  end // always @(posedge)
  assign _cacheEntryMemA_ext_R0_addr = io_in_addr[5:3];
  assign _cacheEntryMemA_ext_W0_en = _GEN_0 | _io_debug_write_T & ~wayReg;
  cacheEntryMem_8x93 cacheEntryMemA_ext (
    .R0_addr (_cacheEntryMemA_ext_R0_addr),
    .R0_en   (_cacheEntryMemA_ext_R0_en),
    .R0_clk  (clock),
    .R0_data (_cacheEntryMemA_ext_R0_data),
    .W0_addr (requestReg_addr_index),
    .W0_en   (_cacheEntryMemA_ext_W0_en),
    .W0_clk  (clock),
    .W0_data (_GEN)
  );
  assign _cacheEntryMemB_ext_R0_addr = io_in_addr[5:3];
  assign _cacheEntryMemB_ext_W0_en = _GEN_0 | _io_debug_write_T & wayReg;
  cacheEntryMem_8x93 cacheEntryMemB_ext (
    .R0_addr (_cacheEntryMemB_ext_R0_addr),
    .R0_en   (_cacheEntryMemB_ext_R0_en),
    .R0_clk  (clock),
    .R0_data (_cacheEntryMemB_ext_R0_data),
    .W0_addr (requestReg_addr_index),
    .W0_en   (_cacheEntryMemB_ext_W0_en),
    .W0_clk  (clock),
    .W0_data (_GEN)
  );
  assign io_in_dout = doutReg;
  assign io_in_wait_n = io_enable & _io_debug_idle_T;
  assign io_in_valid = validReg;
  assign io_out_rd = stateReg == 3'h3;
  assign io_out_addr =
    {requestReg_addr_tag[18:0], requestReg_addr_index, requestReg_addr_offset, 1'h0};
endmodule

