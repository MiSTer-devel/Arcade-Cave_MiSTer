module RegisterFile_1(
  input         clock,
  input         io_mem_wr,
  input  [2:0]  io_mem_addr,
  input  [1:0]  io_mem_mask,
  input  [15:0] io_mem_din,
  output [15:0] io_regs_0,
  output [15:0] io_regs_1,
  output [15:0] io_regs_2,
  output [15:0] io_regs_3,
  output [15:0] io_regs_4,
  output [15:0] io_regs_5
);

  reg  [15:0] regs_0;
  reg  [15:0] regs_1;
  reg  [15:0] regs_2;
  reg  [15:0] regs_3;
  reg  [15:0] regs_4;
  reg  [15:0] regs_5;
  reg  [15:0] regs_6;
  reg  [15:0] regs_7;
  reg  [15:0] casez_tmp;
  always @(*) begin
    casez (io_mem_addr)
      3'b000:
        casez_tmp = regs_0;
      3'b001:
        casez_tmp = regs_1;
      3'b010:
        casez_tmp = regs_2;
      3'b011:
        casez_tmp = regs_3;
      3'b100:
        casez_tmp = regs_4;
      3'b101:
        casez_tmp = regs_5;
      3'b110:
        casez_tmp = regs_6;
      default:
        casez_tmp = regs_7;
    endcase
  end // always @(*)
  wire [7:0]  bytes_1 = io_mem_wr & io_mem_mask[1] ? io_mem_din[15:8] : casez_tmp[15:8];
  wire [7:0]  bytes_0 = io_mem_wr & io_mem_mask[0] ? io_mem_din[7:0] : casez_tmp[7:0];
  wire [15:0] _regs_T = {bytes_1, bytes_0};
  always @(posedge clock) begin
    if (io_mem_addr == 3'h0)
      regs_0 <= _regs_T;
    if (io_mem_addr == 3'h1)
      regs_1 <= _regs_T;
    if (io_mem_addr == 3'h2)
      regs_2 <= _regs_T;
    if (io_mem_addr == 3'h3)
      regs_3 <= _regs_T;
    if (io_mem_addr == 3'h4)
      regs_4 <= _regs_T;
    if (io_mem_addr == 3'h5)
      regs_5 <= _regs_T;
    if (io_mem_addr == 3'h6)
      regs_6 <= _regs_T;
    if (&io_mem_addr)
      regs_7 <= _regs_T;
  end // always @(posedge)
  assign io_regs_0 = regs_0;
  assign io_regs_1 = regs_1;
  assign io_regs_2 = regs_2;
  assign io_regs_3 = regs_3;
  assign io_regs_4 = regs_4;
  assign io_regs_5 = regs_5;
endmodule

