module ChannelController(
  input         clock,
  input         reset,
  input  [7:0]  io_regs_0_pitch,
  input         io_regs_0_flags_keyOn,
  input         io_regs_0_flags_loop,
  input  [7:0]  io_regs_0_level,
  input  [3:0]  io_regs_0_pan,
  input  [23:0] io_regs_0_startAddr,
  input  [23:0] io_regs_0_loopStartAddr,
  input  [23:0] io_regs_0_loopEndAddr,
  input  [23:0] io_regs_0_endAddr,
  input  [7:0]  io_regs_1_pitch,
  input         io_regs_1_flags_keyOn,
  input         io_regs_1_flags_loop,
  input  [7:0]  io_regs_1_level,
  input  [3:0]  io_regs_1_pan,
  input  [23:0] io_regs_1_startAddr,
  input  [23:0] io_regs_1_loopStartAddr,
  input  [23:0] io_regs_1_loopEndAddr,
  input  [23:0] io_regs_1_endAddr,
  input  [7:0]  io_regs_2_pitch,
  input         io_regs_2_flags_keyOn,
  input         io_regs_2_flags_loop,
  input  [7:0]  io_regs_2_level,
  input  [3:0]  io_regs_2_pan,
  input  [23:0] io_regs_2_startAddr,
  input  [23:0] io_regs_2_loopStartAddr,
  input  [23:0] io_regs_2_loopEndAddr,
  input  [23:0] io_regs_2_endAddr,
  input  [7:0]  io_regs_3_pitch,
  input         io_regs_3_flags_keyOn,
  input         io_regs_3_flags_loop,
  input  [7:0]  io_regs_3_level,
  input  [3:0]  io_regs_3_pan,
  input  [23:0] io_regs_3_startAddr,
  input  [23:0] io_regs_3_loopStartAddr,
  input  [23:0] io_regs_3_loopEndAddr,
  input  [23:0] io_regs_3_endAddr,
  input  [7:0]  io_regs_4_pitch,
  input         io_regs_4_flags_keyOn,
  input         io_regs_4_flags_loop,
  input  [7:0]  io_regs_4_level,
  input  [3:0]  io_regs_4_pan,
  input  [23:0] io_regs_4_startAddr,
  input  [23:0] io_regs_4_loopStartAddr,
  input  [23:0] io_regs_4_loopEndAddr,
  input  [23:0] io_regs_4_endAddr,
  input  [7:0]  io_regs_5_pitch,
  input         io_regs_5_flags_keyOn,
  input         io_regs_5_flags_loop,
  input  [7:0]  io_regs_5_level,
  input  [3:0]  io_regs_5_pan,
  input  [23:0] io_regs_5_startAddr,
  input  [23:0] io_regs_5_loopStartAddr,
  input  [23:0] io_regs_5_loopEndAddr,
  input  [23:0] io_regs_5_endAddr,
  input  [7:0]  io_regs_6_pitch,
  input         io_regs_6_flags_keyOn,
  input         io_regs_6_flags_loop,
  input  [7:0]  io_regs_6_level,
  input  [3:0]  io_regs_6_pan,
  input  [23:0] io_regs_6_startAddr,
  input  [23:0] io_regs_6_loopStartAddr,
  input  [23:0] io_regs_6_loopEndAddr,
  input  [23:0] io_regs_6_endAddr,
  input  [7:0]  io_regs_7_pitch,
  input         io_regs_7_flags_keyOn,
  input         io_regs_7_flags_loop,
  input  [7:0]  io_regs_7_level,
  input  [3:0]  io_regs_7_pan,
  input  [23:0] io_regs_7_startAddr,
  input  [23:0] io_regs_7_loopStartAddr,
  input  [23:0] io_regs_7_loopEndAddr,
  input  [23:0] io_regs_7_endAddr,
  input         io_enable,
  output        io_done,
  output [2:0]  io_index,
  output        io_audio_valid,
  output [15:0] io_audio_bits_left,
  output        io_rom_rd,
  output [23:0] io_rom_addr,
  input  [7:0]  io_rom_dout,
  input         io_rom_wait_n,
  input         io_rom_valid
);

  wire         _audioPipeline_io_in_ready;
  wire         _audioPipeline_io_out_valid;
  wire [15:0]  _audioPipeline_io_out_bits_state_samples_0;
  wire [15:0]  _audioPipeline_io_out_bits_state_samples_1;
  wire         _audioPipeline_io_out_bits_state_underflow;
  wire [15:0]  _audioPipeline_io_out_bits_state_adpcmStep;
  wire [9:0]   _audioPipeline_io_out_bits_state_lerpIndex;
  wire         _audioPipeline_io_out_bits_state_loopEnable;
  wire [15:0]  _audioPipeline_io_out_bits_state_loopStep;
  wire [15:0]  _audioPipeline_io_out_bits_state_loopSample;
  wire [16:0]  _audioPipeline_io_out_bits_audio_left;
  wire         _audioPipeline_io_pcmData_ready;
  wire         _channelStateMem_ext_W0_en;
  wire [120:0] _channelStateMem_ext_W0_data;
  wire [120:0] _channelStateMem_ext_R0_data;
  reg  [3:0]   stateReg;
  reg  [16:0]  accumulatorReg_left;
  wire         _io_debug_init_T = stateReg == 4'h0;
  reg  [2:0]   channelCounter;
  reg  [8:0]   outputCounterWrap_value;
  wire         outputCounterWrap = outputCounterWrap_value == 9'h16A;
  wire         _io_debug_read_T = stateReg == 4'h2;
  reg          channelStateReg_enable;
  reg          channelStateReg_active;
  reg          channelStateReg_done;
  reg          channelStateReg_nibble;
  reg  [23:0]  channelStateReg_addr;
  reg          channelStateReg_loopStart;
  reg  [15:0]  channelStateReg_audioPipelineState_samples_0;
  reg  [15:0]  channelStateReg_audioPipelineState_samples_1;
  reg          channelStateReg_audioPipelineState_underflow;
  reg  [15:0]  channelStateReg_audioPipelineState_adpcmStep;
  reg  [9:0]   channelStateReg_audioPipelineState_lerpIndex;
  reg          channelStateReg_audioPipelineState_loopEnable;
  reg  [15:0]  channelStateReg_audioPipelineState_loopStep;
  reg  [15:0]  channelStateReg_audioPipelineState_loopSample;
  wire         audioPipeline_io_in_valid = stateReg == 4'h5;
  reg  [7:0]   casez_tmp;
  always @(*) begin
    casez (channelCounter)
      3'b000:
        casez_tmp = io_regs_0_pitch;
      3'b001:
        casez_tmp = io_regs_1_pitch;
      3'b010:
        casez_tmp = io_regs_2_pitch;
      3'b011:
        casez_tmp = io_regs_3_pitch;
      3'b100:
        casez_tmp = io_regs_4_pitch;
      3'b101:
        casez_tmp = io_regs_5_pitch;
      3'b110:
        casez_tmp = io_regs_6_pitch;
      default:
        casez_tmp = io_regs_7_pitch;
    endcase
  end // always @(*)
  reg          casez_tmp_0;
  always @(*) begin
    casez (channelCounter)
      3'b000:
        casez_tmp_0 = io_regs_0_flags_keyOn;
      3'b001:
        casez_tmp_0 = io_regs_1_flags_keyOn;
      3'b010:
        casez_tmp_0 = io_regs_2_flags_keyOn;
      3'b011:
        casez_tmp_0 = io_regs_3_flags_keyOn;
      3'b100:
        casez_tmp_0 = io_regs_4_flags_keyOn;
      3'b101:
        casez_tmp_0 = io_regs_5_flags_keyOn;
      3'b110:
        casez_tmp_0 = io_regs_6_flags_keyOn;
      default:
        casez_tmp_0 = io_regs_7_flags_keyOn;
    endcase
  end // always @(*)
  reg          casez_tmp_1;
  always @(*) begin
    casez (channelCounter)
      3'b000:
        casez_tmp_1 = io_regs_0_flags_loop;
      3'b001:
        casez_tmp_1 = io_regs_1_flags_loop;
      3'b010:
        casez_tmp_1 = io_regs_2_flags_loop;
      3'b011:
        casez_tmp_1 = io_regs_3_flags_loop;
      3'b100:
        casez_tmp_1 = io_regs_4_flags_loop;
      3'b101:
        casez_tmp_1 = io_regs_5_flags_loop;
      3'b110:
        casez_tmp_1 = io_regs_6_flags_loop;
      default:
        casez_tmp_1 = io_regs_7_flags_loop;
    endcase
  end // always @(*)
  reg  [7:0]   casez_tmp_2;
  always @(*) begin
    casez (channelCounter)
      3'b000:
        casez_tmp_2 = io_regs_0_level;
      3'b001:
        casez_tmp_2 = io_regs_1_level;
      3'b010:
        casez_tmp_2 = io_regs_2_level;
      3'b011:
        casez_tmp_2 = io_regs_3_level;
      3'b100:
        casez_tmp_2 = io_regs_4_level;
      3'b101:
        casez_tmp_2 = io_regs_5_level;
      3'b110:
        casez_tmp_2 = io_regs_6_level;
      default:
        casez_tmp_2 = io_regs_7_level;
    endcase
  end // always @(*)
  reg  [3:0]   casez_tmp_3;
  always @(*) begin
    casez (channelCounter)
      3'b000:
        casez_tmp_3 = io_regs_0_pan;
      3'b001:
        casez_tmp_3 = io_regs_1_pan;
      3'b010:
        casez_tmp_3 = io_regs_2_pan;
      3'b011:
        casez_tmp_3 = io_regs_3_pan;
      3'b100:
        casez_tmp_3 = io_regs_4_pan;
      3'b101:
        casez_tmp_3 = io_regs_5_pan;
      3'b110:
        casez_tmp_3 = io_regs_6_pan;
      default:
        casez_tmp_3 = io_regs_7_pan;
    endcase
  end // always @(*)
  reg  [23:0]  casez_tmp_4;
  always @(*) begin
    casez (channelCounter)
      3'b000:
        casez_tmp_4 = io_regs_0_startAddr;
      3'b001:
        casez_tmp_4 = io_regs_1_startAddr;
      3'b010:
        casez_tmp_4 = io_regs_2_startAddr;
      3'b011:
        casez_tmp_4 = io_regs_3_startAddr;
      3'b100:
        casez_tmp_4 = io_regs_4_startAddr;
      3'b101:
        casez_tmp_4 = io_regs_5_startAddr;
      3'b110:
        casez_tmp_4 = io_regs_6_startAddr;
      default:
        casez_tmp_4 = io_regs_7_startAddr;
    endcase
  end // always @(*)
  reg  [23:0]  casez_tmp_5;
  always @(*) begin
    casez (channelCounter)
      3'b000:
        casez_tmp_5 = io_regs_0_loopStartAddr;
      3'b001:
        casez_tmp_5 = io_regs_1_loopStartAddr;
      3'b010:
        casez_tmp_5 = io_regs_2_loopStartAddr;
      3'b011:
        casez_tmp_5 = io_regs_3_loopStartAddr;
      3'b100:
        casez_tmp_5 = io_regs_4_loopStartAddr;
      3'b101:
        casez_tmp_5 = io_regs_5_loopStartAddr;
      3'b110:
        casez_tmp_5 = io_regs_6_loopStartAddr;
      default:
        casez_tmp_5 = io_regs_7_loopStartAddr;
    endcase
  end // always @(*)
  reg  [23:0]  casez_tmp_6;
  always @(*) begin
    casez (channelCounter)
      3'b000:
        casez_tmp_6 = io_regs_0_loopEndAddr;
      3'b001:
        casez_tmp_6 = io_regs_1_loopEndAddr;
      3'b010:
        casez_tmp_6 = io_regs_2_loopEndAddr;
      3'b011:
        casez_tmp_6 = io_regs_3_loopEndAddr;
      3'b100:
        casez_tmp_6 = io_regs_4_loopEndAddr;
      3'b101:
        casez_tmp_6 = io_regs_5_loopEndAddr;
      3'b110:
        casez_tmp_6 = io_regs_6_loopEndAddr;
      default:
        casez_tmp_6 = io_regs_7_loopEndAddr;
    endcase
  end // always @(*)
  reg  [23:0]  casez_tmp_7;
  always @(*) begin
    casez (channelCounter)
      3'b000:
        casez_tmp_7 = io_regs_0_endAddr;
      3'b001:
        casez_tmp_7 = io_regs_1_endAddr;
      3'b010:
        casez_tmp_7 = io_regs_2_endAddr;
      3'b011:
        casez_tmp_7 = io_regs_3_endAddr;
      3'b100:
        casez_tmp_7 = io_regs_4_endAddr;
      3'b101:
        casez_tmp_7 = io_regs_5_endAddr;
      3'b110:
        casez_tmp_7 = io_regs_6_endAddr;
      default:
        casez_tmp_7 = io_regs_7_endAddr;
    endcase
  end // always @(*)
  wire [3:0]   audioPipeline_io_pcmData_bits =
    channelStateReg_nibble ? io_rom_dout[3:0] : io_rom_dout[7:4];
  reg          pendingReg;
  wire         _io_debug_check_T = stateReg == 4'h4;
  wire         _io_debug_write_T = stateReg == 4'h7;
  wire [23:0]  data_addr = _io_debug_write_T ? channelStateReg_addr : 24'h0;
  wire [15:0]  data_audioPipelineState_samples_0 =
    _io_debug_write_T ? channelStateReg_audioPipelineState_samples_0 : 16'h0;
  wire [15:0]  data_audioPipelineState_samples_1 =
    _io_debug_write_T ? channelStateReg_audioPipelineState_samples_1 : 16'h0;
  wire [15:0]  data_audioPipelineState_adpcmStep =
    _io_debug_write_T ? channelStateReg_audioPipelineState_adpcmStep : 16'h7F;
  wire [9:0]   data_audioPipelineState_lerpIndex =
    _io_debug_write_T ? channelStateReg_audioPipelineState_lerpIndex : 10'h0;
  wire [15:0]  data_audioPipelineState_loopStep =
    _io_debug_write_T ? channelStateReg_audioPipelineState_loopStep : 16'h0;
  wire [15:0]  data_audioPipelineState_loopSample =
    _io_debug_write_T ? channelStateReg_audioPipelineState_loopSample : 16'h0;
  wire [16:0]  _io_audio_bits_T_1 =
    $signed(accumulatorReg_left) < -17'sh8000 ? 17'h18000 : accumulatorReg_left;
  wire         _io_debug_next_T = stateReg == 4'h8;
  wire         _GEN = _io_debug_init_T | _io_debug_next_T;
  wire         channelCounterWrap = _GEN & (&channelCounter);
  wire         _io_debug_latch_T = stateReg == 4'h3;
  wire         _GEN_0 =
    _io_debug_latch_T ? _channelStateMem_ext_R0_data[119] : channelStateReg_active;
  wire         start = ~channelStateReg_enable & ~channelStateReg_active & casez_tmp_0;
  wire         stop = channelStateReg_enable & ~casez_tmp_0;
  wire         _io_debug_idle_T = stateReg == 4'h1;
  wire         _GEN_1 = _io_debug_check_T & start;
  wire         _GEN_2 = _audioPipeline_io_pcmData_ready & io_rom_valid;
  wire         _GEN_3 = casez_tmp_1 & channelStateReg_addr == casez_tmp_6;
  wire         _GEN_4 = channelStateReg_addr == casez_tmp_7;
  wire         _GEN_5 = _GEN_2 & channelStateReg_nibble;
  wire         _GEN_6 =
    _io_debug_latch_T ? _channelStateMem_ext_R0_data[120] : channelStateReg_enable;
  wire         _GEN_7 = _io_debug_check_T ? start | ~stop & _GEN_0 : _GEN_0;
  wire         _GEN_8 =
    _io_debug_latch_T ? _channelStateMem_ext_R0_data[118] : channelStateReg_done;
  wire         _GEN_9 =
    _io_debug_latch_T ? _channelStateMem_ext_R0_data[117] : channelStateReg_nibble;
  wire         _GEN_10 =
    _io_debug_latch_T ? _channelStateMem_ext_R0_data[92] : channelStateReg_loopStart;
  wire         _GEN_11 =
    _io_debug_latch_T
      ? _channelStateMem_ext_R0_data[59]
      : channelStateReg_audioPipelineState_underflow;
  wire         _GEN_12 =
    _io_debug_latch_T
      ? _channelStateMem_ext_R0_data[32]
      : channelStateReg_audioPipelineState_loopEnable;
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 4'h0;
      channelCounter <= 3'h0;
      outputCounterWrap_value <= 9'h0;
      pendingReg <= 1'h0;
    end
    else begin
      if (_io_debug_init_T) begin
        if (channelCounterWrap)
          stateReg <= 4'h1;
      end
      else if (_io_debug_idle_T) begin
        if (io_enable)
          stateReg <= 4'h2;
      end
      else if (_io_debug_read_T)
        stateReg <= 4'h3;
      else if (_io_debug_latch_T)
        stateReg <= 4'h4;
      else if (_io_debug_check_T)
        stateReg <= {2'h1, ~(channelStateReg_active | start), 1'h1};
      else if (audioPipeline_io_in_valid) begin
        if (_audioPipeline_io_in_ready)
          stateReg <= 4'h6;
      end
      else if (stateReg == 4'h6) begin
        if (_audioPipeline_io_out_valid)
          stateReg <= 4'h7;
      end
      else if (_io_debug_write_T)
        stateReg <= 4'h8;
      else if (_io_debug_next_T)
        stateReg <= channelCounterWrap ? 4'h9 : 4'h2;
      else if (stateReg == 4'h9 & outputCounterWrap)
        stateReg <= 4'h1;
      if (_GEN)
        channelCounter <= 3'(channelCounter + 3'h1);
      outputCounterWrap_value <=
        outputCounterWrap ? 9'h0 : 9'(outputCounterWrap_value + 9'h1);
      pendingReg <=
        ~io_rom_valid & (_audioPipeline_io_pcmData_ready & io_rom_wait_n | pendingReg);
    end
    if (_audioPipeline_io_out_valid) begin
      accumulatorReg_left <=
        17'(accumulatorReg_left + _audioPipeline_io_out_bits_audio_left);
      channelStateReg_audioPipelineState_samples_0 <=
        _audioPipeline_io_out_bits_state_samples_0;
      channelStateReg_audioPipelineState_samples_1 <=
        _audioPipeline_io_out_bits_state_samples_1;
      channelStateReg_audioPipelineState_adpcmStep <=
        _audioPipeline_io_out_bits_state_adpcmStep;
      channelStateReg_audioPipelineState_lerpIndex <=
        _audioPipeline_io_out_bits_state_lerpIndex;
      channelStateReg_audioPipelineState_loopStep <=
        _audioPipeline_io_out_bits_state_loopStep;
      channelStateReg_audioPipelineState_loopSample <=
        _audioPipeline_io_out_bits_state_loopSample;
    end
    else begin
      if (_io_debug_idle_T)
        accumulatorReg_left <= 17'h0;
      if (_GEN_1) begin
        channelStateReg_audioPipelineState_samples_0 <= 16'h0;
        channelStateReg_audioPipelineState_samples_1 <= 16'h0;
        channelStateReg_audioPipelineState_adpcmStep <= 16'h7F;
        channelStateReg_audioPipelineState_lerpIndex <= 10'h0;
        channelStateReg_audioPipelineState_loopStep <= 16'h0;
        channelStateReg_audioPipelineState_loopSample <= 16'h0;
      end
      else if (_io_debug_latch_T) begin
        channelStateReg_audioPipelineState_samples_0 <=
          _channelStateMem_ext_R0_data[75:60];
        channelStateReg_audioPipelineState_samples_1 <=
          _channelStateMem_ext_R0_data[91:76];
        channelStateReg_audioPipelineState_adpcmStep <=
          _channelStateMem_ext_R0_data[58:43];
        channelStateReg_audioPipelineState_lerpIndex <=
          _channelStateMem_ext_R0_data[42:33];
        channelStateReg_audioPipelineState_loopStep <=
          _channelStateMem_ext_R0_data[31:16];
        channelStateReg_audioPipelineState_loopSample <=
          _channelStateMem_ext_R0_data[15:0];
      end
    end
    if (_io_debug_check_T)
      channelStateReg_enable <= start | ~stop & _GEN_6;
    else if (_io_debug_latch_T)
      channelStateReg_enable <= _channelStateMem_ext_R0_data[120];
    channelStateReg_active <= (~_GEN_5 | _GEN_3 | ~_GEN_4) & _GEN_7;
    channelStateReg_done <=
      _GEN_5 & ~_GEN_3 & _GEN_4
      | ~(_io_debug_check_T & (start | stop | channelStateReg_done)) & _GEN_8;
    channelStateReg_nibble <= _GEN_2 ? ~channelStateReg_nibble : ~_GEN_1 & _GEN_9;
    if (_GEN_5) begin
      if (_GEN_3)
        channelStateReg_addr <= casez_tmp_5;
      else if (_GEN_4) begin
        if (_GEN_1)
          channelStateReg_addr <= casez_tmp_4;
        else if (_io_debug_latch_T)
          channelStateReg_addr <= _channelStateMem_ext_R0_data[116:93];
      end
      else
        channelStateReg_addr <= 24'(channelStateReg_addr + 24'h1);
    end
    else if (_GEN_1)
      channelStateReg_addr <= casez_tmp_4;
    else if (_io_debug_latch_T)
      channelStateReg_addr <= _channelStateMem_ext_R0_data[116:93];
    channelStateReg_loopStart <=
      _GEN_2
        ? casez_tmp_1 & channelStateReg_addr == casez_tmp_5 & ~channelStateReg_nibble
        : ~_GEN_1 & _GEN_10;
    channelStateReg_audioPipelineState_underflow <=
      _audioPipeline_io_out_valid
        ? _audioPipeline_io_out_bits_state_underflow
        : _GEN_1 | _GEN_11;
    channelStateReg_audioPipelineState_loopEnable <=
      _audioPipeline_io_out_valid
        ? _audioPipeline_io_out_bits_state_loopEnable
        : ~_GEN_1 & _GEN_12;
  end // always @(posedge)
  assign _channelStateMem_ext_W0_en = _io_debug_init_T | _io_debug_write_T;
  assign _channelStateMem_ext_W0_data =
    {_io_debug_write_T & channelStateReg_enable,
     _io_debug_write_T & channelStateReg_active,
     _io_debug_write_T & channelStateReg_done,
     _io_debug_write_T & channelStateReg_nibble,
     data_addr,
     _io_debug_write_T & channelStateReg_loopStart,
     data_audioPipelineState_samples_1,
     data_audioPipelineState_samples_0,
     ~_io_debug_write_T | channelStateReg_audioPipelineState_underflow,
     data_audioPipelineState_adpcmStep,
     data_audioPipelineState_lerpIndex,
     _io_debug_write_T & channelStateReg_audioPipelineState_loopEnable,
     data_audioPipelineState_loopStep,
     data_audioPipelineState_loopSample};
  channelStateMem_8x121 channelStateMem_ext (
    .R0_addr (channelCounter),
    .R0_en   (_io_debug_read_T),
    .R0_clk  (clock),
    .R0_data (_channelStateMem_ext_R0_data),
    .W0_addr (channelCounter),
    .W0_en   (_channelStateMem_ext_W0_en),
    .W0_clk  (clock),
    .W0_data (_channelStateMem_ext_W0_data)
  );
  AudioPipeline audioPipeline (
    .clock                        (clock),
    .reset                        (reset),
    .io_in_ready                  (_audioPipeline_io_in_ready),
    .io_in_valid                  (audioPipeline_io_in_valid),
    .io_in_bits_state_samples_0   (channelStateReg_audioPipelineState_samples_0),
    .io_in_bits_state_samples_1   (channelStateReg_audioPipelineState_samples_1),
    .io_in_bits_state_underflow   (channelStateReg_audioPipelineState_underflow),
    .io_in_bits_state_adpcmStep   (channelStateReg_audioPipelineState_adpcmStep),
    .io_in_bits_state_lerpIndex   (channelStateReg_audioPipelineState_lerpIndex),
    .io_in_bits_state_loopEnable  (channelStateReg_audioPipelineState_loopEnable),
    .io_in_bits_state_loopStep    (channelStateReg_audioPipelineState_loopStep),
    .io_in_bits_state_loopSample  (channelStateReg_audioPipelineState_loopSample),
    .io_in_bits_pitch             (casez_tmp),
    .io_in_bits_level             (casez_tmp_2),
    .io_in_bits_pan               (casez_tmp_3),
    .io_out_valid                 (_audioPipeline_io_out_valid),
    .io_out_bits_state_samples_0  (_audioPipeline_io_out_bits_state_samples_0),
    .io_out_bits_state_samples_1  (_audioPipeline_io_out_bits_state_samples_1),
    .io_out_bits_state_underflow  (_audioPipeline_io_out_bits_state_underflow),
    .io_out_bits_state_adpcmStep  (_audioPipeline_io_out_bits_state_adpcmStep),
    .io_out_bits_state_lerpIndex  (_audioPipeline_io_out_bits_state_lerpIndex),
    .io_out_bits_state_loopEnable (_audioPipeline_io_out_bits_state_loopEnable),
    .io_out_bits_state_loopStep   (_audioPipeline_io_out_bits_state_loopStep),
    .io_out_bits_state_loopSample (_audioPipeline_io_out_bits_state_loopSample),
    .io_out_bits_audio_left       (_audioPipeline_io_out_bits_audio_left),
    .io_pcmData_ready             (_audioPipeline_io_pcmData_ready),
    .io_pcmData_valid             (io_rom_valid),
    .io_pcmData_bits              (audioPipeline_io_pcmData_bits),
    .io_loopStart                 (channelStateReg_loopStart)
  );
  assign io_done = _io_debug_check_T & channelStateReg_done;
  assign io_index = channelCounter;
  assign io_audio_valid = outputCounterWrap;
  assign io_audio_bits_left =
    $signed(_io_audio_bits_T_1) < 17'sh7FFF ? _io_audio_bits_T_1[15:0] : 16'h7FFF;
  assign io_rom_rd = _audioPipeline_io_pcmData_ready & ~pendingReg;
  assign io_rom_addr = channelStateReg_addr;
endmodule

