module Main(
  input   clock,
  input   reset
);
endmodule
