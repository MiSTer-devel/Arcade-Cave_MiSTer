module SpriteFrameBuffer(
  input         clock,
  input         reset,
  input         io_videoClock,
  input         io_enable,
  input         io_swap,
  input  [8:0]  io_video_pos_y,
  input         io_video_hBlank,
  input  [8:0]  io_lineBuffer_addr,
  output [15:0] io_lineBuffer_dout,
  input         io_frameBuffer_wr,
  input  [16:0] io_frameBuffer_addr,
  input  [15:0] io_frameBuffer_din,
  output        io_frameBuffer_wait_n,
  output        io_ddr_rd,
  output        io_ddr_wr,
  output [31:0] io_ddr_addr,
  output [7:0]  io_ddr_mask,
  output [63:0] io_ddr_din,
  input  [63:0] io_ddr_dout,
  input         io_ddr_wait_n,
  input         io_ddr_valid,
  output [7:0]  io_ddr_burstLength,
  input         io_ddr_burstDone
);

  wire [31:0] _ddrArbiter_io_in_0_addr;
  wire [31:0] _ddrArbiter_io_in_1_addr;
  wire [31:0] _ddrArbiter_io_in_2_addr;
  wire        _frameBufferDma_io_out_wait_n;
  wire        _frameBufferDma_io_out_burstDone;
  wire        _frameBufferDma_io_out_wr;
  wire [31:0] _frameBufferDma_io_out_addr;
  wire [63:0] _frameBufferDma_io_out_din;
  wire        _queue_io_out_wait_n;
  wire        _queue_io_out_wr;
  wire [31:0] _queue_io_out_addr;
  wire [7:0]  _queue_io_out_mask;
  wire [63:0] _queue_io_out_din;
  wire        _lineBufferDma_io_start;
  wire [63:0] _lineBufferDma_io_in_dout;
  wire        _lineBufferDma_io_in_wait_n;
  wire        _lineBufferDma_io_in_valid;
  wire        _lineBufferDma_io_in_burstDone;
  wire        _lineBufferDma_io_in_rd;
  wire [31:0] _lineBufferDma_io_in_addr;
  wire [31:0] _lineBufferDma_io_out_addr;
  wire [31:0] _pageFlipper_io_addrRead;
  wire [31:0] _pageFlipper_io_addrWrite;
  wire        _lineBuffer_io_portA_wr;
  wire [6:0]  _lineBuffer_io_portA_addr;
  wire [63:0] _lineBuffer_io_portA_din;
  reg         hBlank_r;
  reg         hBlank;
  reg         hBlankRising_REG;
  wire        frameBufferDma_io_start = io_enable & io_swap;
  always @(posedge clock) begin
    hBlank_r <= io_video_hBlank;
    hBlank <= hBlank_r;
    hBlankRising_REG <= hBlank;
  end // always @(posedge)
  assign _lineBuffer_io_portA_addr = _lineBufferDma_io_out_addr[9:3];
  TrueDualPortRam_11 lineBuffer (
    .clock         (clock),
    .io_clockB     (io_videoClock),
    .io_portA_wr   (_lineBuffer_io_portA_wr),
    .io_portA_addr (_lineBuffer_io_portA_addr),
    .io_portA_din  (_lineBuffer_io_portA_din),
    .io_portB_addr (io_lineBuffer_addr),
    .io_portB_dout (io_lineBuffer_dout)
  );
  PageFlipper pageFlipper (
    .clock        (clock),
    .reset        (reset),
    .io_swapWrite (frameBufferDma_io_start),
    .io_addrRead  (_pageFlipper_io_addrRead),
    .io_addrWrite (_pageFlipper_io_addrWrite)
  );
  assign _lineBufferDma_io_start = io_enable & hBlank & ~hBlankRising_REG;
  BurstReadDMA_1 lineBufferDma (
    .clock           (clock),
    .reset           (reset),
    .io_start        (_lineBufferDma_io_start),
    .io_in_rd        (_lineBufferDma_io_in_rd),
    .io_in_addr      (_lineBufferDma_io_in_addr),
    .io_in_dout      (_lineBufferDma_io_in_dout),
    .io_in_wait_n    (_lineBufferDma_io_in_wait_n),
    .io_in_valid     (_lineBufferDma_io_in_valid),
    .io_in_burstDone (_lineBufferDma_io_in_burstDone),
    .io_out_wr       (_lineBuffer_io_portA_wr),
    .io_out_addr     (_lineBufferDma_io_out_addr),
    .io_out_din      (_lineBuffer_io_portA_din)
  );
  RequestQueue queue (
    .clock         (clock),
    .io_enable     (io_enable),
    .io_readClock  (clock),
    .io_in_wr      (io_frameBuffer_wr),
    .io_in_addr    (io_frameBuffer_addr),
    .io_in_din     (io_frameBuffer_din),
    .io_in_wait_n  (io_frameBuffer_wait_n),
    .io_out_wr     (_queue_io_out_wr),
    .io_out_addr   (_queue_io_out_addr),
    .io_out_mask   (_queue_io_out_mask),
    .io_out_din    (_queue_io_out_din),
    .io_out_wait_n (_queue_io_out_wait_n)
  );
  BurstWriteDMA frameBufferDma (
    .clock            (clock),
    .reset            (reset),
    .io_start         (frameBufferDma_io_start),
    .io_out_wr        (_frameBufferDma_io_out_wr),
    .io_out_addr      (_frameBufferDma_io_out_addr),
    .io_out_din       (_frameBufferDma_io_out_din),
    .io_out_wait_n    (_frameBufferDma_io_out_wait_n),
    .io_out_burstDone (_frameBufferDma_io_out_burstDone)
  );
  assign _ddrArbiter_io_in_0_addr =
    32'(_lineBufferDma_io_in_addr
        + 32'(_pageFlipper_io_addrRead + {13'h0, 9'(io_video_pos_y + 9'h1), 10'h0}));
  assign _ddrArbiter_io_in_1_addr =
    32'(_frameBufferDma_io_out_addr + _pageFlipper_io_addrWrite);
  assign _ddrArbiter_io_in_2_addr = 32'(_queue_io_out_addr + _pageFlipper_io_addrWrite);
  BurstMemArbiter_2 ddrArbiter (
    .clock              (clock),
    .reset              (reset),
    .io_in_0_rd         (_lineBufferDma_io_in_rd),
    .io_in_0_addr       (_ddrArbiter_io_in_0_addr),
    .io_in_0_dout       (_lineBufferDma_io_in_dout),
    .io_in_0_wait_n     (_lineBufferDma_io_in_wait_n),
    .io_in_0_valid      (_lineBufferDma_io_in_valid),
    .io_in_0_burstDone  (_lineBufferDma_io_in_burstDone),
    .io_in_1_wr         (_frameBufferDma_io_out_wr),
    .io_in_1_addr       (_ddrArbiter_io_in_1_addr),
    .io_in_1_din        (_frameBufferDma_io_out_din),
    .io_in_1_wait_n     (_frameBufferDma_io_out_wait_n),
    .io_in_1_burstDone  (_frameBufferDma_io_out_burstDone),
    .io_in_2_wr         (_queue_io_out_wr),
    .io_in_2_addr       (_ddrArbiter_io_in_2_addr),
    .io_in_2_mask       (_queue_io_out_mask),
    .io_in_2_din        (_queue_io_out_din),
    .io_in_2_wait_n     (_queue_io_out_wait_n),
    .io_out_rd          (io_ddr_rd),
    .io_out_wr          (io_ddr_wr),
    .io_out_addr        (io_ddr_addr),
    .io_out_mask        (io_ddr_mask),
    .io_out_din         (io_ddr_din),
    .io_out_dout        (io_ddr_dout),
    .io_out_wait_n      (io_ddr_wait_n),
    .io_out_valid       (io_ddr_valid),
    .io_out_burstLength (io_ddr_burstLength),
    .io_out_burstDone   (io_ddr_burstDone)
  );
endmodule

