module RegisterFile(
  input         clock,
  input         io_mem_wr,
  input  [1:0]  io_mem_addr,
  input  [15:0] io_mem_din,
  output [15:0] io_regs_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] regs_0; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_1; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_2; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_3; // @[RegisterFile.scala 56:17]
  wire [15:0] _GEN_1 = 2'h1 == io_mem_addr ? regs_1 : regs_0; // @[]
  wire [15:0] _GEN_2 = 2'h2 == io_mem_addr ? regs_2 : _GEN_1; // @[]
  wire [15:0] _GEN_3 = 2'h3 == io_mem_addr ? regs_3 : _GEN_2; // @[]
  wire [7:0] bytes_0 = io_mem_wr ? io_mem_din[7:0] : _GEN_3[7:0]; // @[RegisterFile.scala 62:28 66:{39,50}]
  wire [7:0] bytes_1 = io_mem_wr ? io_mem_din[15:8] : _GEN_3[15:8]; // @[RegisterFile.scala 62:28 66:{39,50}]
  wire [15:0] _regs_T = {bytes_1,bytes_0}; // @[RegisterFile.scala 70:17]
  assign io_regs_0 = regs_0; // @[RegisterFile.scala 74:11]
  always @(posedge clock) begin
    if (2'h0 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_0 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (2'h1 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_1 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (2'h2 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_2 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (2'h3 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_3 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DDR(
  input         clock,
  input         reset,
  input         io_mem_rd,
  input         io_mem_wr,
  input  [31:0] io_mem_addr,
  input  [7:0]  io_mem_mask,
  input  [63:0] io_mem_din,
  output [63:0] io_mem_dout,
  output        io_mem_wait_n,
  output        io_mem_valid,
  input  [7:0]  io_mem_burstLength,
  output        io_mem_burstDone,
  output        io_ddr_rd,
  output        io_ddr_wr,
  output [31:0] io_ddr_addr,
  output [7:0]  io_ddr_mask,
  output [63:0] io_ddr_din,
  input  [63:0] io_ddr_dout,
  input         io_ddr_wait_n,
  input         io_ddr_valid,
  output [7:0]  io_ddr_burstLength
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[DDR.scala 62:25]
  wire  _burstLength_T = stateReg == 2'h0; // @[DDR.scala 63:34]
  reg [7:0] burstLength_r; // @[Reg.scala 19:16]
  wire [7:0] _GEN_0 = _burstLength_T ? io_mem_burstLength : burstLength_r; // @[Reg.scala 19:16 20:{18,22}]
  wire  read = _burstLength_T & io_mem_rd; // @[DDR.scala 69:38]
  wire  write = (_burstLength_T | stateReg == 2'h2) & io_mem_wr; // @[DDR.scala 70:73]
  wire  effectiveRead = read & io_ddr_wait_n; // @[DDR.scala 71:28]
  wire  effectiveWrite = write & io_ddr_wait_n; // @[DDR.scala 72:30]
  wire  burstCounterEnable = stateReg == 2'h1 & io_ddr_valid | effectiveWrite; // @[DDR.scala 73:74]
  reg [7:0] burstCounter; // @[Counter.scala 65:22]
  wire [7:0] _wrap_wrap_T_1 = _GEN_0 - 8'h1; // @[Counter.scala 69:29]
  wire  wrap_wrap = burstCounter == _wrap_wrap_T_1 | _GEN_0 == 8'h0; // @[Counter.scala 69:35]
  wire [7:0] _wrap_value_T_1 = burstCounter + 8'h1; // @[Counter.scala 70:20]
  wire  burstCounterWrap = burstCounterEnable & wrap_wrap; // @[Counter.scala 93:{48,55}]
  assign io_mem_dout = io_ddr_dout; // @[DDR.scala 86:10]
  assign io_mem_wait_n = io_ddr_wait_n; // @[DDR.scala 86:10]
  assign io_mem_valid = io_ddr_valid; // @[DDR.scala 86:10]
  assign io_mem_burstDone = burstCounterEnable & wrap_wrap; // @[Counter.scala 93:{48,55}]
  assign io_ddr_rd = _burstLength_T & io_mem_rd; // @[DDR.scala 69:38]
  assign io_ddr_wr = (_burstLength_T | stateReg == 2'h2) & io_mem_wr; // @[DDR.scala 70:73]
  assign io_ddr_addr = io_mem_addr; // @[DDR.scala 86:10]
  assign io_ddr_mask = io_mem_mask; // @[DDR.scala 86:10]
  assign io_ddr_din = io_mem_din; // @[DDR.scala 86:10]
  assign io_ddr_burstLength = stateReg == 2'h0 ? io_mem_burstLength : burstLength_r; // @[DDR.scala 63:24]
  always @(posedge clock) begin
    if (reset) begin // @[DDR.scala 62:25]
      stateReg <= 2'h0; // @[DDR.scala 62:25]
    end else if (burstCounterWrap) begin // @[Mux.scala 101:16]
      stateReg <= 2'h0;
    end else if (effectiveRead) begin // @[Mux.scala 101:16]
      stateReg <= 2'h1;
    end else if (effectiveWrite) begin // @[Mux.scala 101:16]
      stateReg <= 2'h2;
    end
    if (_burstLength_T) begin // @[Reg.scala 20:18]
      burstLength_r <= io_mem_burstLength; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[Counter.scala 65:22]
      burstCounter <= 8'h0; // @[Counter.scala 65:22]
    end else if (burstCounterEnable) begin // @[Counter.scala 93:48]
      if (wrap_wrap) begin // @[Counter.scala 71:16]
        burstCounter <= 8'h0; // @[Counter.scala 71:24]
      end else begin
        burstCounter <= _wrap_value_T_1; // @[Counter.scala 70:11]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  burstLength_r = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  burstCounter = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SDRAM(
  input         clock,
  input         reset,
  input         io_mem_rd,
  input         io_mem_wr,
  input  [24:0] io_mem_addr,
  input  [15:0] io_mem_din,
  output [15:0] io_mem_dout,
  output        io_mem_wait_n,
  output        io_mem_valid,
  output        io_mem_burstDone,
  output        io_sdram_cs_n,
  output        io_sdram_ras_n,
  output        io_sdram_cas_n,
  output        io_sdram_we_n,
  output        io_sdram_oe_n,
  output [1:0]  io_sdram_bank,
  output [12:0] io_sdram_addr,
  output [15:0] io_sdram_din,
  input  [15:0] io_sdram_dout
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] stateReg; // @[SDRAM.scala 79:25]
  reg [3:0] commandReg; // @[SDRAM.scala 83:27]
  reg [14:0] waitCounter; // @[Counter.scala 40:34]
  wire  _T_1 = waitCounter == 15'h0; // @[SDRAM.scala 186:24]
  wire [2:0] _GEN_16 = waitCounter == 15'h4b0d ? 3'h1 : stateReg; // @[SDRAM.scala 194:128 140:13 147:15]
  wire [2:0] _GEN_19 = waitCounter == 15'h4b07 ? stateReg : _GEN_16; // @[SDRAM.scala 192:107 140:13]
  wire [2:0] _GEN_22 = waitCounter == 15'h4b01 ? stateReg : _GEN_19; // @[SDRAM.scala 140:13 190:86]
  wire [2:0] _GEN_25 = waitCounter == 15'h4aff ? stateReg : _GEN_22; // @[SDRAM.scala 140:13 188:63]
  wire [2:0] _GEN_28 = waitCounter == 15'h0 ? stateReg : _GEN_25; // @[SDRAM.scala 140:13 186:33]
  wire  modeDone = waitCounter == 15'h1; // @[SDRAM.scala 112:30]
  wire [2:0] _GEN_30 = modeDone ? 3'h2 : stateReg; // @[SDRAM.scala 140:13 152:15 201:22]
  reg [9:0] refreshCounter; // @[Counter.scala 40:34]
  wire  triggerRefresh = refreshCounter >= 10'h2eb; // @[SDRAM.scala 117:39]
  wire  isReadWrite = io_mem_rd | io_mem_wr; // @[SDRAM.scala 89:31]
  wire [2:0] _GEN_32 = isReadWrite ? 3'h3 : stateReg; // @[SDRAM.scala 140:13 157:15 206:64]
  wire [2:0] _GEN_36 = triggerRefresh ? 3'h6 : _GEN_32; // @[SDRAM.scala 178:15 206:28]
  reg  requestReg_wr; // @[Reg.scala 19:16]
  wire [2:0] _GEN_40 = requestReg_wr ? 3'h5 : 3'h4; // @[SDRAM.scala 164:15 171:15 212:29]
  wire [2:0] _GEN_44 = modeDone ? _GEN_40 : stateReg; // @[SDRAM.scala 140:13 211:24]
  wire  readDone = waitCounter == 15'h5; // @[SDRAM.scala 114:30]
  wire [2:0] _GEN_47 = isReadWrite ? 3'h3 : 3'h2; // @[SDRAM.scala 152:15 157:15 219:66]
  wire [2:0] _GEN_48 = triggerRefresh ? 3'h6 : _GEN_47; // @[SDRAM.scala 178:15 219:30]
  wire [2:0] _GEN_50 = readDone ? _GEN_48 : stateReg; // @[SDRAM.scala 140:13 218:22]
  wire  writeDone = waitCounter == 15'h6; // @[SDRAM.scala 115:31]
  wire [2:0] _GEN_54 = writeDone ? _GEN_48 : stateReg; // @[SDRAM.scala 140:13 225:23]
  wire [2:0] _GEN_58 = readDone ? _GEN_47 : stateReg; // @[SDRAM.scala 140:13 232:25]
  wire [2:0] _GEN_62 = 3'h6 == stateReg ? _GEN_58 : stateReg; // @[SDRAM.scala 140:13 182:20]
  wire [2:0] _GEN_66 = 3'h5 == stateReg ? _GEN_54 : _GEN_62; // @[SDRAM.scala 182:20]
  wire [2:0] _GEN_70 = 3'h4 == stateReg ? _GEN_50 : _GEN_66; // @[SDRAM.scala 182:20]
  wire [2:0] _GEN_74 = 3'h3 == stateReg ? _GEN_44 : _GEN_70; // @[SDRAM.scala 182:20]
  wire [2:0] _GEN_78 = 3'h2 == stateReg ? _GEN_36 : _GEN_74; // @[SDRAM.scala 182:20]
  wire [2:0] _GEN_81 = 3'h1 == stateReg ? _GEN_30 : _GEN_78; // @[SDRAM.scala 182:20]
  wire [2:0] nextState = 3'h0 == stateReg ? _GEN_28 : _GEN_81; // @[SDRAM.scala 182:20]
  wire  latch = stateReg != 3'h3 & nextState == 3'h3; // @[SDRAM.scala 86:41]
  wire [8:0] request_addr_col = io_mem_addr[9:1]; // @[Address.scala 57:25]
  wire [12:0] request_addr_row = io_mem_addr[22:10]; // @[Address.scala 57:25]
  wire [1:0] request_addr_bank = io_mem_addr[24:23]; // @[Address.scala 57:25]
  reg [1:0] requestReg_addr_bank; // @[Reg.scala 19:16]
  reg [8:0] requestReg_addr_col; // @[Reg.scala 19:16]
  reg [1:0] bankReg; // @[SDRAM.scala 99:20]
  reg [12:0] addrReg; // @[SDRAM.scala 100:20]
  reg [15:0] dinReg; // @[SDRAM.scala 101:23]
  reg [15:0] doutReg; // @[SDRAM.scala 102:24]
  wire  waitCounter_x2 = nextState != stateReg; // @[SDRAM.scala 105:82]
  wire [14:0] _waitCounter_wrap_value_T_1 = waitCounter + 15'h1; // @[Counter.scala 46:22]
  wire  _refreshCounter_T_2 = stateReg != 3'h0 & stateReg != 3'h1; // @[SDRAM.scala 107:38]
  wire  _refreshCounter_T_5 = stateReg == 3'h6 & _T_1; // @[SDRAM.scala 108:40]
  wire [9:0] _refreshCounter_wrap_value_T_1 = refreshCounter + 10'h1; // @[Counter.scala 46:22]
  wire  burstBusy = waitCounter < 15'h3; // @[SDRAM.scala 118:31]
  wire  burstDone = waitCounter == 15'h3; // @[SDRAM.scala 119:31]
  wire  wait_n_idle = stateReg == 3'h2 & ~isReadWrite; // @[SDRAM.scala 123:40]
  wire  wait_n_read = latch & io_mem_rd; // @[SDRAM.scala 124:22]
  wire  _wait_n_write_T_3 = stateReg == 3'h5; // @[SDRAM.scala 125:89]
  wire  wait_n_write = stateReg == 3'h3 & modeDone & requestReg_wr | stateReg == 3'h5 & burstBusy; // @[SDRAM.scala 125:76]
  wire  _validReg_T = stateReg == 3'h4; // @[SDRAM.scala 130:35]
  reg  validReg; // @[SDRAM.scala 130:25]
  wire  memBurstDone_readBurstDone = _validReg_T & readDone; // @[SDRAM.scala 134:49]
  wire  memBurstDone_writeBurstDone = _wait_n_write_T_3 & burstDone; // @[SDRAM.scala 135:51]
  reg  memBurstDone_REG; // @[SDRAM.scala 136:12]
  wire [3:0] _GEN_15 = waitCounter == 15'h4b0d ? 4'h0 : 4'h7; // @[SDRAM.scala 194:128 143:15 146:17]
  wire [12:0] _GEN_17 = waitCounter == 15'h4b0d ? 13'h22 : 13'h400; // @[SDRAM.scala 194:128 148:13 185:15]
  wire [3:0] _GEN_18 = waitCounter == 15'h4b07 ? 4'h1 : _GEN_15; // @[SDRAM.scala 192:107 193:21]
  wire [12:0] _GEN_20 = waitCounter == 15'h4b07 ? 13'h400 : _GEN_17; // @[SDRAM.scala 192:107 185:15]
  wire [3:0] _GEN_21 = waitCounter == 15'h4b01 ? 4'h1 : _GEN_18; // @[SDRAM.scala 190:86 191:21]
  wire [3:0] _GEN_31 = isReadWrite ? 4'h3 : 4'h7; // @[SDRAM.scala 143:15 156:17 206:64]
  wire [1:0] _GEN_33 = isReadWrite ? request_addr_bank : bankReg; // @[SDRAM.scala 158:13 206:64 99:20]
  wire [12:0] _GEN_34 = isReadWrite ? request_addr_row : addrReg; // @[SDRAM.scala 159:13 100:20 206:64]
  wire [3:0] _GEN_35 = triggerRefresh ? 4'h1 : _GEN_31; // @[SDRAM.scala 177:17 206:28]
  wire [1:0] _GEN_37 = triggerRefresh ? bankReg : _GEN_33; // @[SDRAM.scala 206:28 99:20]
  wire [12:0] _GEN_38 = triggerRefresh ? addrReg : _GEN_34; // @[SDRAM.scala 100:20 206:28]
  wire [9:0] _addrReg_T_5 = {{1'd0}, requestReg_addr_col}; // @[SDRAM.scala 173:51]
  wire [10:0] _addrReg_T_6 = {1'h1,_addrReg_T_5}; // @[SDRAM.scala 173:25]
  wire [3:0] _GEN_39 = requestReg_wr ? 4'h4 : 4'h5; // @[SDRAM.scala 163:17 170:17 212:29]
  wire [10:0] _GEN_42 = requestReg_wr ? _addrReg_T_6 : _addrReg_T_6; // @[SDRAM.scala 166:13 173:13 212:29]
  wire [3:0] _GEN_43 = modeDone ? _GEN_39 : 4'h7; // @[SDRAM.scala 143:15 211:24]
  wire [1:0] _GEN_45 = modeDone ? requestReg_addr_bank : bankReg; // @[SDRAM.scala 211:24 99:20]
  wire [12:0] _GEN_46 = modeDone ? {{2'd0}, _GEN_42} : addrReg; // @[SDRAM.scala 100:20 211:24]
  wire [3:0] _GEN_49 = readDone ? _GEN_35 : 4'h7; // @[SDRAM.scala 143:15 218:22]
  wire [1:0] _GEN_51 = readDone ? _GEN_37 : bankReg; // @[SDRAM.scala 218:22 99:20]
  wire [12:0] _GEN_52 = readDone ? _GEN_38 : addrReg; // @[SDRAM.scala 100:20 218:22]
  wire [3:0] _GEN_53 = writeDone ? _GEN_35 : 4'h7; // @[SDRAM.scala 143:15 225:23]
  wire [1:0] _GEN_55 = writeDone ? _GEN_37 : bankReg; // @[SDRAM.scala 225:23 99:20]
  wire [12:0] _GEN_56 = writeDone ? _GEN_38 : addrReg; // @[SDRAM.scala 100:20 225:23]
  wire [3:0] _GEN_57 = readDone ? _GEN_31 : 4'h7; // @[SDRAM.scala 143:15 232:25]
  wire [1:0] _GEN_59 = readDone ? _GEN_33 : bankReg; // @[SDRAM.scala 232:25 99:20]
  wire [12:0] _GEN_60 = readDone ? _GEN_34 : addrReg; // @[SDRAM.scala 100:20 232:25]
  wire [3:0] _GEN_61 = 3'h6 == stateReg ? _GEN_57 : 4'h7; // @[SDRAM.scala 143:15 182:20]
  wire [1:0] _GEN_63 = 3'h6 == stateReg ? _GEN_59 : bankReg; // @[SDRAM.scala 182:20 99:20]
  wire [12:0] _GEN_64 = 3'h6 == stateReg ? _GEN_60 : addrReg; // @[SDRAM.scala 100:20 182:20]
  wire [3:0] _GEN_65 = 3'h5 == stateReg ? _GEN_53 : _GEN_61; // @[SDRAM.scala 182:20]
  wire [1:0] _GEN_67 = 3'h5 == stateReg ? _GEN_55 : _GEN_63; // @[SDRAM.scala 182:20]
  wire [12:0] _GEN_68 = 3'h5 == stateReg ? _GEN_56 : _GEN_64; // @[SDRAM.scala 182:20]
  wire [3:0] _GEN_69 = 3'h4 == stateReg ? _GEN_49 : _GEN_65; // @[SDRAM.scala 182:20]
  wire [1:0] _GEN_71 = 3'h4 == stateReg ? _GEN_51 : _GEN_67; // @[SDRAM.scala 182:20]
  wire [12:0] _GEN_72 = 3'h4 == stateReg ? _GEN_52 : _GEN_68; // @[SDRAM.scala 182:20]
  wire [3:0] _GEN_73 = 3'h3 == stateReg ? _GEN_43 : _GEN_69; // @[SDRAM.scala 182:20]
  assign io_mem_dout = doutReg; // @[SDRAM.scala 242:15]
  assign io_mem_wait_n = wait_n_idle | wait_n_read | wait_n_write; // @[SDRAM.scala 126:18]
  assign io_mem_valid = validReg; // @[SDRAM.scala 240:16]
  assign io_mem_burstDone = memBurstDone_REG | memBurstDone_writeBurstDone; // @[SDRAM.scala 136:37]
  assign io_sdram_cs_n = commandReg[3]; // @[SDRAM.scala 244:30]
  assign io_sdram_ras_n = commandReg[2]; // @[SDRAM.scala 245:31]
  assign io_sdram_cas_n = commandReg[1]; // @[SDRAM.scala 246:31]
  assign io_sdram_we_n = commandReg[0]; // @[SDRAM.scala 247:30]
  assign io_sdram_oe_n = stateReg != 3'h4; // @[SDRAM.scala 248:29]
  assign io_sdram_bank = bankReg; // @[SDRAM.scala 249:17]
  assign io_sdram_addr = addrReg; // @[SDRAM.scala 250:17]
  assign io_sdram_din = dinReg; // @[SDRAM.scala 251:16]
  always @(posedge clock) begin
    if (reset) begin // @[SDRAM.scala 79:25]
      stateReg <= 3'h0; // @[SDRAM.scala 79:25]
    end else if (3'h0 == stateReg) begin // @[SDRAM.scala 182:20]
      if (!(waitCounter == 15'h0)) begin // @[SDRAM.scala 186:33]
        if (!(waitCounter == 15'h4aff)) begin // @[SDRAM.scala 188:63]
          stateReg <= _GEN_22;
        end
      end
    end else if (3'h1 == stateReg) begin // @[SDRAM.scala 182:20]
      if (modeDone) begin // @[SDRAM.scala 201:22]
        stateReg <= 3'h2; // @[SDRAM.scala 152:15]
      end
    end else if (3'h2 == stateReg) begin // @[SDRAM.scala 182:20]
      stateReg <= _GEN_36;
    end else begin
      stateReg <= _GEN_74;
    end
    if (reset) begin // @[SDRAM.scala 83:27]
      commandReg <= 4'h7; // @[SDRAM.scala 83:27]
    end else if (3'h0 == stateReg) begin // @[SDRAM.scala 182:20]
      if (waitCounter == 15'h0) begin // @[SDRAM.scala 186:33]
        commandReg <= 4'h8; // @[SDRAM.scala 187:21]
      end else if (waitCounter == 15'h4aff) begin // @[SDRAM.scala 188:63]
        commandReg <= 4'h2; // @[SDRAM.scala 189:21]
      end else begin
        commandReg <= _GEN_21;
      end
    end else if (3'h1 == stateReg) begin // @[SDRAM.scala 182:20]
      commandReg <= 4'h7; // @[SDRAM.scala 143:15]
    end else if (3'h2 == stateReg) begin // @[SDRAM.scala 182:20]
      commandReg <= _GEN_35;
    end else begin
      commandReg <= _GEN_73;
    end
    if (reset) begin // @[Counter.scala 40:34]
      waitCounter <= 15'h0; // @[Counter.scala 40:34]
    end else if (waitCounter_x2) begin // @[Counter.scala 86:17]
      waitCounter <= 15'h0; // @[Counter.scala 59:13]
    end else begin
      waitCounter <= _waitCounter_wrap_value_T_1;
    end
    if (reset) begin // @[Counter.scala 40:34]
      refreshCounter <= 10'h0; // @[Counter.scala 40:34]
    end else if (_refreshCounter_T_5) begin // @[Counter.scala 86:17]
      refreshCounter <= 10'h0; // @[Counter.scala 59:13]
    end else if (_refreshCounter_T_2) begin // @[Counter.scala 86:48]
      refreshCounter <= _refreshCounter_wrap_value_T_1; // @[Counter.scala 46:13]
    end
    if (latch) begin // @[Reg.scala 20:18]
      requestReg_wr <= io_mem_wr; // @[Reg.scala 20:22]
    end
    if (latch) begin // @[Reg.scala 20:18]
      requestReg_addr_bank <= request_addr_bank; // @[Reg.scala 20:22]
    end
    if (latch) begin // @[Reg.scala 20:18]
      requestReg_addr_col <= request_addr_col; // @[Reg.scala 20:22]
    end
    if (!(3'h0 == stateReg)) begin // @[SDRAM.scala 182:20]
      if (!(3'h1 == stateReg)) begin // @[SDRAM.scala 182:20]
        if (3'h2 == stateReg) begin // @[SDRAM.scala 182:20]
          if (!(triggerRefresh)) begin // @[SDRAM.scala 206:28]
            bankReg <= _GEN_33;
          end
        end else if (3'h3 == stateReg) begin // @[SDRAM.scala 182:20]
          bankReg <= _GEN_45;
        end else begin
          bankReg <= _GEN_71;
        end
      end
    end
    if (3'h0 == stateReg) begin // @[SDRAM.scala 182:20]
      if (waitCounter == 15'h0) begin // @[SDRAM.scala 186:33]
        addrReg <= 13'h400; // @[SDRAM.scala 185:15]
      end else if (waitCounter == 15'h4aff) begin // @[SDRAM.scala 188:63]
        addrReg <= 13'h400; // @[SDRAM.scala 185:15]
      end else if (waitCounter == 15'h4b01) begin // @[SDRAM.scala 190:86]
        addrReg <= 13'h400; // @[SDRAM.scala 185:15]
      end else begin
        addrReg <= _GEN_20;
      end
    end else if (!(3'h1 == stateReg)) begin // @[SDRAM.scala 182:20]
      if (3'h2 == stateReg) begin // @[SDRAM.scala 182:20]
        if (!(triggerRefresh)) begin // @[SDRAM.scala 206:28]
          addrReg <= _GEN_34;
        end
      end else if (3'h3 == stateReg) begin // @[SDRAM.scala 182:20]
        addrReg <= _GEN_46;
      end else begin
        addrReg <= _GEN_72;
      end
    end
    dinReg <= io_mem_din; // @[SDRAM.scala 101:23]
    doutReg <= io_sdram_dout; // @[SDRAM.scala 102:24]
    if (reset) begin // @[SDRAM.scala 130:25]
      validReg <= 1'h0; // @[SDRAM.scala 130:25]
    end else begin
      validReg <= stateReg == 3'h4 & waitCounter > 15'h1; // @[SDRAM.scala 130:25]
    end
    if (reset) begin // @[SDRAM.scala 136:12]
      memBurstDone_REG <= 1'h0; // @[SDRAM.scala 136:12]
    end else begin
      memBurstDone_REG <= memBurstDone_readBurstDone; // @[SDRAM.scala 136:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  commandReg = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  waitCounter = _RAND_2[14:0];
  _RAND_3 = {1{`RANDOM}};
  refreshCounter = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  requestReg_wr = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  requestReg_addr_bank = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  requestReg_addr_col = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  bankReg = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  addrReg = _RAND_8[12:0];
  _RAND_9 = {1{`RANDOM}};
  dinReg = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  doutReg = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  validReg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  memBurstDone_REG = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BurstBuffer(
  input         clock,
  input         reset,
  input         io_in_wr,
  input  [26:0] io_in_addr,
  input  [15:0] io_in_din,
  output        io_out_wr,
  output [31:0] io_out_addr,
  output [63:0] io_out_din,
  input         io_out_burstDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  writePendingReg; // @[BurstBuffer.scala 56:32]
  reg [63:0] lineReg_words_0; // @[BurstBuffer.scala 57:20]
  reg [26:0] addrReg; // @[BurstBuffer.scala 58:20]
  reg  busyReg; // @[BurstBuffer.scala 59:24]
  wire  latchAddr = io_in_wr & ~busyReg; // @[BurstBuffer.scala 62:28]
  wire  latchData = io_in_wr & ~writePendingReg; // @[BurstBuffer.scala 63:28]
  reg [1:0] wordCounter; // @[Counter.scala 40:34]
  wire  wrap_wrap = wordCounter == 2'h3; // @[Counter.scala 45:24]
  wire [1:0] _wrap_value_T_1 = wordCounter + 2'h1; // @[Counter.scala 46:22]
  wire  wordCounterWrap = latchData & wrap_wrap; // @[Counter.scala 86:{48,55}]
  wire  _GEN_6 = io_in_wr | busyReg; // @[BurstBuffer.scala 73:24 74:13 59:24]
  wire  _GEN_8 = wordCounterWrap | writePendingReg; // @[BurstBuffer.scala 80:31 81:21 56:32]
  wire [15:0] words_ws_0 = lineReg_words_0[15:0]; // @[Util.scala 104:11]
  wire [15:0] words_ws_1 = lineReg_words_0[31:16]; // @[Util.scala 104:11]
  wire [15:0] words_ws_2 = lineReg_words_0[47:32]; // @[Util.scala 104:11]
  wire [15:0] words_ws_3 = lineReg_words_0[63:48]; // @[Util.scala 104:11]
  wire [15:0] words_0 = 2'h0 == wordCounter ? io_in_din : words_ws_0; // @[BurstBuffer.scala 92:{24,24}]
  wire [15:0] words_1 = 2'h1 == wordCounter ? io_in_din : words_ws_1; // @[BurstBuffer.scala 92:{24,24}]
  wire [15:0] words_2 = 2'h2 == wordCounter ? io_in_din : words_ws_2; // @[BurstBuffer.scala 92:{24,24}]
  wire [15:0] words_3 = 2'h3 == wordCounter ? io_in_din : words_ws_3; // @[BurstBuffer.scala 92:{24,24}]
  wire [63:0] _T = {words_3,words_2,words_1,words_0}; // @[BurstBuffer.scala 93:36]
  wire [26:0] _io_out_addr_T_1 = {addrReg[26:3], 3'h0}; // @[Util.scala 135:64]
  assign io_out_wr = writePendingReg; // @[BurstBuffer.scala 98:13]
  assign io_out_addr = {{5'd0}, _io_out_addr_T_1}; // @[BurstBuffer.scala 100:15]
  assign io_out_din = lineReg_words_0; // @[BurstBuffer.scala 101:14]
  always @(posedge clock) begin
    if (reset) begin // @[BurstBuffer.scala 56:32]
      writePendingReg <= 1'h0; // @[BurstBuffer.scala 56:32]
    end else if (io_out_burstDone) begin // @[BurstBuffer.scala 78:26]
      writePendingReg <= 1'h0; // @[BurstBuffer.scala 79:21]
    end else begin
      writePendingReg <= _GEN_8;
    end
    if (latchData) begin // @[BurstBuffer.scala 90:19]
      lineReg_words_0 <= _T; // @[BurstBuffer.scala 93:19]
    end
    if (latchAddr) begin // @[BurstBuffer.scala 85:19]
      addrReg <= io_in_addr; // @[BurstBuffer.scala 86:13]
    end
    if (reset) begin // @[BurstBuffer.scala 59:24]
      busyReg <= 1'h0; // @[BurstBuffer.scala 59:24]
    end else if (io_out_burstDone) begin // @[BurstBuffer.scala 71:26]
      busyReg <= 1'h0; // @[BurstBuffer.scala 72:13]
    end else begin
      busyReg <= _GEN_6;
    end
    if (reset) begin // @[Counter.scala 40:34]
      wordCounter <= 2'h0; // @[Counter.scala 40:34]
    end else if (latchData) begin // @[Counter.scala 86:48]
      wordCounter <= _wrap_value_T_1; // @[Counter.scala 46:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writePendingReg = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  lineReg_words_0 = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  addrReg = _RAND_2[26:0];
  _RAND_3 = {1{`RANDOM}};
  busyReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wordCounter = _RAND_4[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BurstBuffer_1(
  input         clock,
  input         reset,
  input         io_in_wr,
  input  [31:0] io_in_addr,
  input  [63:0] io_in_din,
  output        io_in_wait_n,
  output        io_out_wr,
  output [24:0] io_out_addr,
  output [15:0] io_out_din,
  input         io_out_wait_n,
  input         io_out_burstDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  writePendingReg; // @[BurstBuffer.scala 56:32]
  reg [15:0] lineReg_words_0; // @[BurstBuffer.scala 57:20]
  reg [15:0] lineReg_words_1; // @[BurstBuffer.scala 57:20]
  reg [15:0] lineReg_words_2; // @[BurstBuffer.scala 57:20]
  reg [15:0] lineReg_words_3; // @[BurstBuffer.scala 57:20]
  reg [31:0] addrReg; // @[BurstBuffer.scala 58:20]
  reg  busyReg; // @[BurstBuffer.scala 59:24]
  wire  latchAddr = io_in_wr & ~busyReg; // @[BurstBuffer.scala 62:28]
  wire  latchData = io_in_wr & ~writePendingReg; // @[BurstBuffer.scala 63:28]
  wire  effectiveWrite = writePendingReg & io_out_wait_n; // @[BurstBuffer.scala 64:40]
  reg [1:0] burstCounter; // @[Counter.scala 40:34]
  wire [1:0] _wrap_value_T_1 = burstCounter + 2'h1; // @[Counter.scala 46:22]
  wire  _GEN_6 = io_in_wr | busyReg; // @[BurstBuffer.scala 73:24 74:13 59:24]
  wire  _GEN_8 = latchData | writePendingReg; // @[BurstBuffer.scala 80:31 81:21 56:32]
  wire [31:0] _io_out_addr_T_1 = {addrReg[31:1], 1'h0}; // @[Util.scala 135:64]
  wire [15:0] _GEN_16 = 2'h1 == burstCounter ? lineReg_words_1 : lineReg_words_0; // @[BurstBuffer.scala 101:{14,14}]
  wire [15:0] _GEN_17 = 2'h2 == burstCounter ? lineReg_words_2 : _GEN_16; // @[BurstBuffer.scala 101:{14,14}]
  assign io_in_wait_n = ~writePendingReg; // @[BurstBuffer.scala 97:19]
  assign io_out_wr = writePendingReg; // @[BurstBuffer.scala 98:13]
  assign io_out_addr = _io_out_addr_T_1[24:0]; // @[BurstBuffer.scala 100:15]
  assign io_out_din = 2'h3 == burstCounter ? lineReg_words_3 : _GEN_17; // @[BurstBuffer.scala 101:{14,14}]
  always @(posedge clock) begin
    if (reset) begin // @[BurstBuffer.scala 56:32]
      writePendingReg <= 1'h0; // @[BurstBuffer.scala 56:32]
    end else if (io_out_burstDone) begin // @[BurstBuffer.scala 78:26]
      writePendingReg <= 1'h0; // @[BurstBuffer.scala 79:21]
    end else begin
      writePendingReg <= _GEN_8;
    end
    if (latchData) begin // @[BurstBuffer.scala 90:19]
      lineReg_words_0 <= io_in_din[15:0]; // @[BurstBuffer.scala 93:19]
    end
    if (latchData) begin // @[BurstBuffer.scala 90:19]
      lineReg_words_1 <= io_in_din[31:16]; // @[BurstBuffer.scala 93:19]
    end
    if (latchData) begin // @[BurstBuffer.scala 90:19]
      lineReg_words_2 <= io_in_din[47:32]; // @[BurstBuffer.scala 93:19]
    end
    if (latchData) begin // @[BurstBuffer.scala 90:19]
      lineReg_words_3 <= io_in_din[63:48]; // @[BurstBuffer.scala 93:19]
    end
    if (latchAddr) begin // @[BurstBuffer.scala 85:19]
      addrReg <= io_in_addr; // @[BurstBuffer.scala 86:13]
    end
    if (reset) begin // @[BurstBuffer.scala 59:24]
      busyReg <= 1'h0; // @[BurstBuffer.scala 59:24]
    end else if (io_out_burstDone) begin // @[BurstBuffer.scala 71:26]
      busyReg <= 1'h0; // @[BurstBuffer.scala 72:13]
    end else begin
      busyReg <= _GEN_6;
    end
    if (reset) begin // @[Counter.scala 40:34]
      burstCounter <= 2'h0; // @[Counter.scala 40:34]
    end else if (effectiveWrite) begin // @[Counter.scala 86:48]
      burstCounter <= _wrap_value_T_1; // @[Counter.scala 46:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writePendingReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  lineReg_words_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  lineReg_words_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  lineReg_words_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  lineReg_words_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  addrReg = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  busyReg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  burstCounter = _RAND_7[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits,
  output [5:0]  io_count,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:31]; // @[Decoupled.scala 275:44]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:44]
  wire [4:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:44]
  wire [63:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:44]
  wire [63:0] ram_MPORT_data; // @[Decoupled.scala 275:44]
  wire [4:0] ram_MPORT_addr; // @[Decoupled.scala 275:44]
  wire  ram_MPORT_mask; // @[Decoupled.scala 275:44]
  wire  ram_MPORT_en; // @[Decoupled.scala 275:44]
  reg  ram_io_deq_bits_MPORT_en_pipe_0;
  reg [4:0] ram_io_deq_bits_MPORT_addr_pipe_0;
  reg [4:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [4:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 278:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 279:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 280:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 281:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  wire [4:0] _value_T_1 = enq_ptr_value + 5'h1; // @[Counter.scala 77:24]
  wire [4:0] _value_T_3 = deq_ptr_value + 5'h1; // @[Counter.scala 77:24]
  wire [5:0] _deq_ptr_next_T_1 = 6'h20 - 6'h1; // @[Decoupled.scala 308:57]
  wire [5:0] _GEN_15 = {{1'd0}, deq_ptr_value}; // @[Decoupled.scala 308:42]
  wire [4:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 328:32]
  wire [5:0] _io_count_T_1 = maybe_full & ptr_match ? 6'h20 : 6'h0; // @[Decoupled.scala 331:20]
  wire [5:0] _GEN_16 = {{1'd0}, ptr_diff}; // @[Decoupled.scala 331:62]
  assign ram_io_deq_bits_MPORT_en = ram_io_deq_bits_MPORT_en_pipe_0;
  assign ram_io_deq_bits_MPORT_addr = ram_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:44]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 305:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 304:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_count = _io_count_T_1 | _GEN_16; // @[Decoupled.scala 331:62]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 275:44]
    end
    ram_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_15 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 308:27]
          ram_io_deq_bits_MPORT_addr_pipe_0 <= 5'h0;
        end else begin
          ram_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 298:15]
      enq_ptr_value <= 5'h0; // @[Counter.scala 98:11]
    end else if (do_enq) begin // @[Decoupled.scala 288:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 298:15]
      deq_ptr_value <= 5'h0; // @[Counter.scala 98:11]
    end else if (do_deq) begin // @[Decoupled.scala 292:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 278:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 278:27]
    end else if (io_flush) begin // @[Decoupled.scala 298:15]
      maybe_full <= 1'h0; // @[Decoupled.scala 301:16]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 295:27]
      maybe_full <= do_enq; // @[Decoupled.scala 296:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_io_deq_bits_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_io_deq_bits_MPORT_addr_pipe_0 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BurstReadDMA(
  input         clock,
  input         reset,
  input         io_start,
  output        io_busy,
  output        io_in_rd,
  output [31:0] io_in_addr,
  input  [63:0] io_in_dout,
  input         io_in_wait_n,
  input         io_in_valid,
  input         io_in_burstDone,
  output        io_out_wr,
  output [31:0] io_out_addr,
  output [63:0] io_out_din,
  input         io_out_wait_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  fifo_clock; // @[BurstReadDMA.scala 69:20]
  wire  fifo_reset; // @[BurstReadDMA.scala 69:20]
  wire  fifo_io_enq_ready; // @[BurstReadDMA.scala 69:20]
  wire  fifo_io_enq_valid; // @[BurstReadDMA.scala 69:20]
  wire [63:0] fifo_io_enq_bits; // @[BurstReadDMA.scala 69:20]
  wire  fifo_io_deq_ready; // @[BurstReadDMA.scala 69:20]
  wire  fifo_io_deq_valid; // @[BurstReadDMA.scala 69:20]
  wire [63:0] fifo_io_deq_bits; // @[BurstReadDMA.scala 69:20]
  wire [5:0] fifo_io_count; // @[BurstReadDMA.scala 69:20]
  wire  fifo_io_flush; // @[BurstReadDMA.scala 69:20]
  reg  readEnableReg; // @[BurstReadDMA.scala 62:30]
  reg  writeEnableReg; // @[BurstReadDMA.scala 63:31]
  reg  readPendingReg; // @[BurstReadDMA.scala 64:31]
  wire  fifoAlmostEmpty = fifo_io_count <= 6'h10; // @[BurstReadDMA.scala 70:39]
  wire  busy = readEnableReg | writeEnableReg; // @[BurstReadDMA.scala 73:28]
  wire  start = io_start & ~busy; // @[BurstReadDMA.scala 74:24]
  wire  read = readEnableReg & ~readPendingReg & fifoAlmostEmpty; // @[BurstReadDMA.scala 75:47]
  wire  write = writeEnableReg & fifo_io_deq_valid; // @[BurstReadDMA.scala 76:30]
  wire  effectiveRead = read & io_in_wait_n; // @[BurstReadDMA.scala 77:28]
  wire  effectiveWrite = write & io_out_wait_n; // @[BurstReadDMA.scala 78:30]
  reg [21:0] wordCounter; // @[Counter.scala 40:34]
  wire  wrap_wrap = wordCounter == 22'h3fffff; // @[Counter.scala 45:24]
  wire [21:0] _wrap_value_T_1 = wordCounter + 22'h1; // @[Counter.scala 46:22]
  wire  wordCounterWrap = effectiveWrite & wrap_wrap; // @[Counter.scala 86:{48,55}]
  reg [17:0] burstCounter; // @[Counter.scala 40:34]
  wire  wrap_wrap_1 = burstCounter == 18'h3ffff; // @[Counter.scala 45:24]
  wire [17:0] _wrap_value_T_3 = burstCounter + 18'h1; // @[Counter.scala 46:22]
  wire  burstCounterWrap = io_in_burstDone & wrap_wrap_1; // @[Counter.scala 86:{48,55}]
  wire [24:0] readAddr = {burstCounter, 7'h0}; // @[BurstReadDMA.scala 87:19]
  wire [24:0] writeAddr = {wordCounter, 3'h0}; // @[BurstReadDMA.scala 93:18]
  wire  _GEN_8 = burstCounterWrap ? 1'h0 : readEnableReg; // @[BurstReadDMA.scala 100:{70,86} 62:30]
  wire  _GEN_9 = start | _GEN_8; // @[BurstReadDMA.scala 100:{15,31}]
  wire  _GEN_10 = wordCounterWrap ? 1'h0 : writeEnableReg; // @[BurstReadDMA.scala 101:{70,87} 63:31]
  wire  _GEN_11 = start | _GEN_10; // @[BurstReadDMA.scala 101:{15,32}]
  wire  _GEN_12 = effectiveRead | readPendingReg; // @[BurstReadDMA.scala 106:29 107:20 64:31]
  Queue fifo ( // @[BurstReadDMA.scala 69:20]
    .clock(fifo_clock),
    .reset(fifo_reset),
    .io_enq_ready(fifo_io_enq_ready),
    .io_enq_valid(fifo_io_enq_valid),
    .io_enq_bits(fifo_io_enq_bits),
    .io_deq_ready(fifo_io_deq_ready),
    .io_deq_valid(fifo_io_deq_valid),
    .io_deq_bits(fifo_io_deq_bits),
    .io_count(fifo_io_count),
    .io_flush(fifo_io_flush)
  );
  assign io_busy = readEnableReg | writeEnableReg; // @[BurstReadDMA.scala 73:28]
  assign io_in_rd = readEnableReg & ~readPendingReg & fifoAlmostEmpty; // @[BurstReadDMA.scala 75:47]
  assign io_in_addr = {{7'd0}, readAddr}; // @[BurstReadDMA.scala 124:14]
  assign io_out_wr = writeEnableReg & fifo_io_deq_valid; // @[BurstReadDMA.scala 76:30]
  assign io_out_addr = {{7'd0}, writeAddr}; // @[BurstReadDMA.scala 126:15]
  assign io_out_din = fifo_io_deq_bits; // @[BurstReadDMA.scala 127:14]
  assign fifo_clock = clock;
  assign fifo_reset = reset;
  assign fifo_io_enq_valid = io_in_valid & readPendingReg; // @[BurstReadDMA.scala 111:20]
  assign fifo_io_enq_bits = io_in_dout; // @[BurstReadDMA.scala 111:39 Decoupled.scala 66:19]
  assign fifo_io_deq_ready = write & io_out_wait_n; // @[BurstReadDMA.scala 78:30]
  assign fifo_io_flush = io_start & ~busy; // @[BurstReadDMA.scala 74:24]
  always @(posedge clock) begin
    if (reset) begin // @[BurstReadDMA.scala 62:30]
      readEnableReg <= 1'h0; // @[BurstReadDMA.scala 62:30]
    end else begin
      readEnableReg <= _GEN_9;
    end
    if (reset) begin // @[BurstReadDMA.scala 63:31]
      writeEnableReg <= 1'h0; // @[BurstReadDMA.scala 63:31]
    end else begin
      writeEnableReg <= _GEN_11;
    end
    if (reset) begin // @[BurstReadDMA.scala 64:31]
      readPendingReg <= 1'h0; // @[BurstReadDMA.scala 64:31]
    end else if (io_in_burstDone) begin // @[BurstReadDMA.scala 104:25]
      readPendingReg <= 1'h0; // @[BurstReadDMA.scala 105:20]
    end else begin
      readPendingReg <= _GEN_12;
    end
    if (reset) begin // @[Counter.scala 40:34]
      wordCounter <= 22'h0; // @[Counter.scala 40:34]
    end else if (effectiveWrite) begin // @[Counter.scala 86:48]
      wordCounter <= _wrap_value_T_1; // @[Counter.scala 46:13]
    end
    if (reset) begin // @[Counter.scala 40:34]
      burstCounter <= 18'h0; // @[Counter.scala 40:34]
    end else if (io_in_burstDone) begin // @[Counter.scala 86:48]
      burstCounter <= _wrap_value_T_3; // @[Counter.scala 46:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  readEnableReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  writeEnableReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  readPendingReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  wordCounter = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  burstCounter = _RAND_4[17:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReadCache(
  input         clock,
  input         reset,
  input         io_enable,
  input         io_in_rd,
  input  [19:0] io_in_addr,
  output [15:0] io_in_dout,
  output        io_in_wait_n,
  output        io_in_valid,
  output        io_out_rd,
  output [24:0] io_out_addr,
  input  [15:0] io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [127:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
`endif // RANDOMIZE_REG_INIT
  reg  cacheEntryMemA_valid [0:127]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [6:0] cacheEntryMemA_valid_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_MPORT_data; // @[ReadCache.scala 112:35]
  wire [6:0] cacheEntryMemA_valid_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_valid_cacheEntryA_en_pipe_0;
  reg [6:0] cacheEntryMemA_valid_cacheEntryA_addr_pipe_0;
  reg [10:0] cacheEntryMemA_tag [0:127]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_tag_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [6:0] cacheEntryMemA_tag_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [10:0] cacheEntryMemA_tag_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [10:0] cacheEntryMemA_tag_MPORT_data; // @[ReadCache.scala 112:35]
  wire [6:0] cacheEntryMemA_tag_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_tag_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_tag_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_tag_cacheEntryA_en_pipe_0;
  reg [6:0] cacheEntryMemA_tag_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_0 [0:127]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_0_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [6:0] cacheEntryMemA_line_words_0_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_0_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_0_MPORT_data; // @[ReadCache.scala 112:35]
  wire [6:0] cacheEntryMemA_line_words_0_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_0_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_0_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0;
  reg [6:0] cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_1 [0:127]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_1_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [6:0] cacheEntryMemA_line_words_1_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_1_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_1_MPORT_data; // @[ReadCache.scala 112:35]
  wire [6:0] cacheEntryMemA_line_words_1_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_1_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_1_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0;
  reg [6:0] cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_2 [0:127]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_2_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [6:0] cacheEntryMemA_line_words_2_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_2_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_2_MPORT_data; // @[ReadCache.scala 112:35]
  wire [6:0] cacheEntryMemA_line_words_2_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_2_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_2_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0;
  reg [6:0] cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_3 [0:127]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_3_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [6:0] cacheEntryMemA_line_words_3_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_3_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_3_MPORT_data; // @[ReadCache.scala 112:35]
  wire [6:0] cacheEntryMemA_line_words_3_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_3_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_3_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0;
  reg [6:0] cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0;
  reg  cacheEntryMemB_valid [0:127]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [6:0] cacheEntryMemB_valid_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [6:0] cacheEntryMemB_valid_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_valid_cacheEntryB_en_pipe_0;
  reg [6:0] cacheEntryMemB_valid_cacheEntryB_addr_pipe_0;
  reg [10:0] cacheEntryMemB_tag [0:127]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_tag_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [6:0] cacheEntryMemB_tag_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [10:0] cacheEntryMemB_tag_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [10:0] cacheEntryMemB_tag_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [6:0] cacheEntryMemB_tag_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_tag_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_tag_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_tag_cacheEntryB_en_pipe_0;
  reg [6:0] cacheEntryMemB_tag_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_0 [0:127]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_0_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [6:0] cacheEntryMemB_line_words_0_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_0_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_0_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [6:0] cacheEntryMemB_line_words_0_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_0_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_0_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0;
  reg [6:0] cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_1 [0:127]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_1_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [6:0] cacheEntryMemB_line_words_1_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_1_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_1_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [6:0] cacheEntryMemB_line_words_1_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_1_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_1_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0;
  reg [6:0] cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_2 [0:127]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_2_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [6:0] cacheEntryMemB_line_words_2_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_2_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_2_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [6:0] cacheEntryMemB_line_words_2_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_2_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_2_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0;
  reg [6:0] cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_3 [0:127]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_3_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [6:0] cacheEntryMemB_line_words_3_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_3_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_3_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [6:0] cacheEntryMemB_line_words_3_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_3_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_3_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0;
  reg [6:0] cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0;
  reg [2:0] stateReg; // @[ReadCache.scala 84:25]
  wire [18:0] offsetReg_addr = io_in_addr[19:1]; // @[ReadCache.scala 91:27]
  wire [1:0] offsetReg_offset = offsetReg_addr[1:0]; // @[ReadCache.scala 92:22]
  reg [1:0] offsetReg; // @[Reg.scala 19:16]
  wire  _start_T_1 = stateReg == 3'h1; // @[ReadCache.scala 142:48]
  wire  start = io_enable & io_in_rd & stateReg == 3'h1; // @[ReadCache.scala 142:36]
  wire [19:0] _request_WIRE_1 = {{1'd0}, offsetReg_addr};
  wire [1:0] request_addr_offset = _request_WIRE_1[1:0]; // @[Address.scala 78:49]
  wire [6:0] request_addr_index = _request_WIRE_1[8:2]; // @[Address.scala 78:49]
  wire [10:0] request_addr_tag = _request_WIRE_1[19:9]; // @[Address.scala 78:49]
  reg  requestReg_rd; // @[Reg.scala 19:16]
  reg [10:0] requestReg_addr_tag; // @[Reg.scala 19:16]
  reg [6:0] requestReg_addr_index; // @[Reg.scala 19:16]
  reg [1:0] requestReg_addr_offset; // @[Reg.scala 19:16]
  reg [15:0] doutReg; // @[ReadCache.scala 101:20]
  reg  validReg; // @[ReadCache.scala 102:25]
  reg [127:0] lruReg; // @[ReadCache.scala 105:19]
  reg  wayReg; // @[ReadCache.scala 109:23]
  wire [127:0] _nextWay_T = lruReg >> request_addr_index; // @[ReadCache.scala 169:31]
  wire  _nextWay_T_2 = start ? _nextWay_T[0] : wayReg; // @[ReadCache.scala 169:17]
  wire  hitA = cacheEntryMemA_valid_cacheEntryA_data & cacheEntryMemA_tag_cacheEntryA_data == requestReg_addr_tag; // @[Entry.scala 59:42]
  wire  hitB = cacheEntryMemB_valid_cacheEntryB_data & cacheEntryMemB_tag_cacheEntryB_data == requestReg_addr_tag; // @[Entry.scala 59:42]
  wire  hit = hitA | hitB; // @[ReadCache.scala 146:18]
  wire  _GEN_76 = hit ? ~hitA : _nextWay_T_2; // @[ReadCache.scala 169:11 185:13 207:17]
  wire  _GEN_86 = 3'h2 == stateReg ? _GEN_76 : _nextWay_T_2; // @[ReadCache.scala 169:11 194:20]
  wire  _GEN_91 = 3'h1 == stateReg ? _nextWay_T_2 : _GEN_86; // @[ReadCache.scala 169:11 194:20]
  wire  nextWay = 3'h0 == stateReg ? _nextWay_T_2 : _GEN_91; // @[ReadCache.scala 169:11 194:20]
  wire  _cacheEntryReg_T_valid = nextWay ? cacheEntryMemB_valid_cacheEntryB_data : cacheEntryMemA_valid_cacheEntryA_data
    ; // @[ReadCache.scala 121:36]
  wire  _cacheEntryReg_T_1 = stateReg == 3'h2; // @[ReadCache.scala 121:82]
  reg  cacheEntryReg_valid; // @[Reg.scala 19:16]
  reg [10:0] cacheEntryReg_tag; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_0; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_1; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_2; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_3; // @[Reg.scala 19:16]
  wire  _GEN_10 = _cacheEntryReg_T_1 ? _cacheEntryReg_T_valid : cacheEntryReg_valid; // @[Reg.scala 19:16 20:{18,22}]
  wire  _nextCacheEntry_T = stateReg == 3'h5; // @[ReadCache.scala 124:37]
  wire  _T = stateReg == 3'h0; // @[ReadCache.scala 126:17]
  wire  _T_2 = ~wayReg; // @[ReadCache.scala 126:64]
  wire  _T_3 = _nextCacheEntry_T & ~wayReg; // @[ReadCache.scala 126:61]
  wire  _T_7 = _nextCacheEntry_T & wayReg; // @[ReadCache.scala 130:61]
  wire  burstCounterEnable = stateReg == 3'h4 & io_out_valid; // @[ReadCache.scala 135:56]
  reg [6:0] initCounter; // @[Counter.scala 61:40]
  wire  wrap_wrap = initCounter == 7'h7f; // @[Counter.scala 73:24]
  wire [6:0] _wrap_value_T_1 = initCounter + 7'h1; // @[Counter.scala 77:24]
  wire  initCounterWrap = _T & wrap_wrap; // @[Counter.scala 118:{16,23}]
  reg [1:0] burstCounter; // @[Counter.scala 61:40]
  wire  wrap_wrap_1 = burstCounter == 2'h3; // @[Counter.scala 73:24]
  wire [1:0] _wrap_value_T_3 = burstCounter + 2'h1; // @[Counter.scala 77:24]
  wire  burstCounterWrap = burstCounterEnable & wrap_wrap_1; // @[Counter.scala 118:{16,23}]
  wire  miss = ~hit; // @[ReadCache.scala 147:14]
  wire  wordDone = burstCounter == 2'h0; // @[ReadCache.scala 153:18]
  wire [19:0] _outAddr_T = {requestReg_addr_tag,requestReg_addr_index,requestReg_addr_offset}; // @[ReadCache.scala 165:11]
  wire [20:0] outAddr = {_outAddr_T, 1'h0}; // @[ReadCache.scala 165:18]
  wire [1:0] n = requestReg_addr_offset + burstCounter; // @[ReadCache.scala 173:57]
  wire [15:0] entry_line_words_0 = 2'h0 == n ? io_out_dout : cacheEntryReg_line_words_0; // @[Entry.scala 92:11 93:{30,30}]
  wire [15:0] entry_line_words_1 = 2'h1 == n ? io_out_dout : cacheEntryReg_line_words_1; // @[Entry.scala 92:11 93:{30,30}]
  wire [15:0] entry_line_words_2 = 2'h2 == n ? io_out_dout : cacheEntryReg_line_words_2; // @[Entry.scala 92:11 93:{30,30}]
  wire [15:0] entry_line_words_3 = 2'h3 == n ? io_out_dout : cacheEntryReg_line_words_3; // @[Entry.scala 92:11 93:{30,30}]
  wire [63:0] _doutReg_ws_T = {entry_line_words_3,entry_line_words_2,entry_line_words_1,entry_line_words_0}; // @[Line.scala 77:32]
  wire [15:0] doutReg_ws_0 = _doutReg_ws_T[15:0]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_1 = _doutReg_ws_T[31:16]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_2 = _doutReg_ws_T[47:32]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_3 = _doutReg_ws_T[63:48]; // @[Util.scala 104:11]
  wire [15:0] _GEN_48 = 2'h1 == offsetReg ? doutReg_ws_1 : doutReg_ws_0; // @[Util.scala 104:{11,11}]
  wire [15:0] _GEN_49 = 2'h2 == offsetReg ? doutReg_ws_2 : _GEN_48; // @[Util.scala 104:{11,11}]
  wire [15:0] _GEN_50 = 2'h3 == offsetReg ? doutReg_ws_3 : _GEN_49; // @[Util.scala 104:{11,11}]
  wire [15:0] _doutReg_T_2 = {_GEN_50[7:0],_GEN_50[15:8]}; // @[Util.scala 114:49]
  wire [15:0] _GEN_58 = burstCounterEnable ? _doutReg_T_2 : doutReg; // @[ReadCache.scala 172:53 176:13 101:20]
  wire  _GEN_59 = burstCounterEnable & (requestReg_rd & wordDone); // @[ReadCache.scala 172:53 177:14 102:25]
  wire [63:0] _doutReg_ws_T_1 = {cacheEntryMemA_line_words_3_cacheEntryA_data,
    cacheEntryMemA_line_words_2_cacheEntryA_data,cacheEntryMemA_line_words_1_cacheEntryA_data,
    cacheEntryMemA_line_words_0_cacheEntryA_data}; // @[Line.scala 77:32]
  wire [15:0] doutReg_ws_0_1 = _doutReg_ws_T_1[15:0]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_1_1 = _doutReg_ws_T_1[31:16]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_2_1 = _doutReg_ws_T_1[47:32]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_3_1 = _doutReg_ws_T_1[63:48]; // @[Util.scala 104:11]
  wire [15:0] _GEN_63 = 2'h1 == offsetReg ? doutReg_ws_1_1 : doutReg_ws_0_1; // @[Util.scala 104:{11,11}]
  wire [15:0] _GEN_64 = 2'h2 == offsetReg ? doutReg_ws_2_1 : _GEN_63; // @[Util.scala 104:{11,11}]
  wire [15:0] _GEN_65 = 2'h3 == offsetReg ? doutReg_ws_3_1 : _GEN_64; // @[Util.scala 104:{11,11}]
  wire [15:0] _doutReg_T_5 = {_GEN_65[7:0],_GEN_65[15:8]}; // @[Util.scala 114:49]
  wire [63:0] _doutReg_ws_T_2 = {cacheEntryMemB_line_words_3_cacheEntryB_data,
    cacheEntryMemB_line_words_2_cacheEntryB_data,cacheEntryMemB_line_words_1_cacheEntryB_data,
    cacheEntryMemB_line_words_0_cacheEntryB_data}; // @[Line.scala 77:32]
  wire [15:0] doutReg_ws_0_2 = _doutReg_ws_T_2[15:0]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_1_2 = _doutReg_ws_T_2[31:16]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_2_2 = _doutReg_ws_T_2[47:32]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_3_2 = _doutReg_ws_T_2[63:48]; // @[Util.scala 104:11]
  wire [15:0] _GEN_67 = 2'h1 == offsetReg ? doutReg_ws_1_2 : doutReg_ws_0_2; // @[Util.scala 104:{11,11}]
  wire [15:0] _GEN_68 = 2'h2 == offsetReg ? doutReg_ws_2_2 : _GEN_67; // @[Util.scala 104:{11,11}]
  wire [15:0] _GEN_69 = 2'h3 == offsetReg ? doutReg_ws_3_2 : _GEN_68; // @[Util.scala 104:{11,11}]
  wire [15:0] _doutReg_T_8 = {_GEN_69[7:0],_GEN_69[15:8]}; // @[Util.scala 114:49]
  wire [15:0] _doutReg_T_9 = hitA ? _doutReg_T_5 : _doutReg_T_8; // @[ReadCache.scala 182:19]
  wire [127:0] _lruReg_T = 128'h1 << requestReg_addr_index; // @[ReadCache.scala 184:28]
  wire [127:0] _lruReg_T_1 = lruReg | _lruReg_T; // @[ReadCache.scala 184:28]
  wire [127:0] _lruReg_T_2 = ~lruReg; // @[ReadCache.scala 184:28]
  wire [127:0] _lruReg_T_3 = _lruReg_T_2 | _lruReg_T; // @[ReadCache.scala 184:28]
  wire [127:0] _lruReg_T_4 = ~_lruReg_T_3; // @[ReadCache.scala 184:28]
  wire [127:0] _lruReg_T_5 = hitA ? _lruReg_T_1 : _lruReg_T_4; // @[ReadCache.scala 184:28]
  wire [127:0] _lruReg_T_12 = _T_2 ? _lruReg_T_1 : _lruReg_T_4; // @[ReadCache.scala 190:28]
  wire [2:0] _GEN_70 = miss ? 3'h3 : stateReg; // @[ReadCache.scala 189:14 207:44 84:25]
  wire [127:0] _GEN_71 = miss ? _lruReg_T_12 : lruReg; // @[ReadCache.scala 190:12 105:19 207:44]
  wire [2:0] _GEN_72 = hit ? 3'h1 : _GEN_70; // @[ReadCache.scala 181:14 207:17]
  wire  _GEN_74 = hit | _GEN_59; // @[ReadCache.scala 183:14 207:17]
  wire [2:0] _GEN_77 = io_out_wait_n ? 3'h4 : stateReg; // @[ReadCache.scala 212:{27,38} 84:25]
  wire [2:0] _GEN_78 = burstCounterWrap ? 3'h5 : stateReg; // @[ReadCache.scala 217:{30,41} 84:25]
  wire [2:0] _GEN_79 = 3'h5 == stateReg ? 3'h1 : stateReg; // @[ReadCache.scala 194:20 221:32 84:25]
  wire [2:0] _GEN_80 = 3'h4 == stateReg ? _GEN_78 : _GEN_79; // @[ReadCache.scala 194:20]
  wire [2:0] _GEN_81 = 3'h3 == stateReg ? _GEN_77 : _GEN_80; // @[ReadCache.scala 194:20]
  assign cacheEntryMemA_valid_cacheEntryA_en = cacheEntryMemA_valid_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_valid_cacheEntryA_addr = cacheEntryMemA_valid_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_valid_cacheEntryA_data = cacheEntryMemA_valid[cacheEntryMemA_valid_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_valid_MPORT_data = _nextCacheEntry_T & cacheEntryReg_valid;
  assign cacheEntryMemA_valid_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_valid_MPORT_mask = 1'h1;
  assign cacheEntryMemA_valid_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_tag_cacheEntryA_en = cacheEntryMemA_tag_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_tag_cacheEntryA_addr = cacheEntryMemA_tag_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_tag_cacheEntryA_data = cacheEntryMemA_tag[cacheEntryMemA_tag_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_tag_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_tag : 11'h0;
  assign cacheEntryMemA_tag_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_tag_MPORT_mask = 1'h1;
  assign cacheEntryMemA_tag_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_0_cacheEntryA_en = cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_0_cacheEntryA_addr = cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_0_cacheEntryA_data =
    cacheEntryMemA_line_words_0[cacheEntryMemA_line_words_0_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_line_words_0_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_0 : 16'h0;
  assign cacheEntryMemA_line_words_0_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_0_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_0_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_1_cacheEntryA_en = cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_1_cacheEntryA_addr = cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_1_cacheEntryA_data =
    cacheEntryMemA_line_words_1[cacheEntryMemA_line_words_1_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_line_words_1_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_1 : 16'h0;
  assign cacheEntryMemA_line_words_1_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_1_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_1_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_2_cacheEntryA_en = cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_2_cacheEntryA_addr = cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_2_cacheEntryA_data =
    cacheEntryMemA_line_words_2[cacheEntryMemA_line_words_2_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_line_words_2_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_2 : 16'h0;
  assign cacheEntryMemA_line_words_2_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_2_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_2_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_3_cacheEntryA_en = cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_3_cacheEntryA_addr = cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_3_cacheEntryA_data =
    cacheEntryMemA_line_words_3[cacheEntryMemA_line_words_3_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_line_words_3_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_3 : 16'h0;
  assign cacheEntryMemA_line_words_3_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_3_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_3_MPORT_en = _T | _T_3;
  assign cacheEntryMemB_valid_cacheEntryB_en = cacheEntryMemB_valid_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_valid_cacheEntryB_addr = cacheEntryMemB_valid_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_valid_cacheEntryB_data = cacheEntryMemB_valid[cacheEntryMemB_valid_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_valid_MPORT_1_data = _nextCacheEntry_T & cacheEntryReg_valid;
  assign cacheEntryMemB_valid_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_valid_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_valid_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_tag_cacheEntryB_en = cacheEntryMemB_tag_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_tag_cacheEntryB_addr = cacheEntryMemB_tag_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_tag_cacheEntryB_data = cacheEntryMemB_tag[cacheEntryMemB_tag_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_tag_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_tag : 11'h0;
  assign cacheEntryMemB_tag_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_tag_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_tag_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_0_cacheEntryB_en = cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_0_cacheEntryB_addr = cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_0_cacheEntryB_data =
    cacheEntryMemB_line_words_0[cacheEntryMemB_line_words_0_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_line_words_0_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_0 : 16'h0;
  assign cacheEntryMemB_line_words_0_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_0_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_0_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_1_cacheEntryB_en = cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_1_cacheEntryB_addr = cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_1_cacheEntryB_data =
    cacheEntryMemB_line_words_1[cacheEntryMemB_line_words_1_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_line_words_1_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_1 : 16'h0;
  assign cacheEntryMemB_line_words_1_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_1_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_1_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_2_cacheEntryB_en = cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_2_cacheEntryB_addr = cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_2_cacheEntryB_data =
    cacheEntryMemB_line_words_2[cacheEntryMemB_line_words_2_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_line_words_2_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_2 : 16'h0;
  assign cacheEntryMemB_line_words_2_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_2_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_2_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_3_cacheEntryB_en = cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_3_cacheEntryB_addr = cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_3_cacheEntryB_data =
    cacheEntryMemB_line_words_3[cacheEntryMemB_line_words_3_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_line_words_3_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_3 : 16'h0;
  assign cacheEntryMemB_line_words_3_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_3_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_3_MPORT_1_en = _T | _T_7;
  assign io_in_dout = doutReg; // @[ReadCache.scala 227:14]
  assign io_in_wait_n = io_enable & _start_T_1; // @[ReadCache.scala 143:26]
  assign io_in_valid = validReg; // @[ReadCache.scala 226:15]
  assign io_out_rd = stateReg == 3'h3; // @[ReadCache.scala 228:25]
  assign io_out_addr = {{4'd0}, outAddr}; // @[ReadCache.scala 230:15]
  always @(posedge clock) begin
    if (cacheEntryMemA_valid_MPORT_en & cacheEntryMemA_valid_MPORT_mask) begin
      cacheEntryMemA_valid[cacheEntryMemA_valid_MPORT_addr] <= cacheEntryMemA_valid_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_valid_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_valid_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[8:2];
    end
    if (cacheEntryMemA_tag_MPORT_en & cacheEntryMemA_tag_MPORT_mask) begin
      cacheEntryMemA_tag[cacheEntryMemA_tag_MPORT_addr] <= cacheEntryMemA_tag_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_tag_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_tag_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[8:2];
    end
    if (cacheEntryMemA_line_words_0_MPORT_en & cacheEntryMemA_line_words_0_MPORT_mask) begin
      cacheEntryMemA_line_words_0[cacheEntryMemA_line_words_0_MPORT_addr] <= cacheEntryMemA_line_words_0_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[8:2];
    end
    if (cacheEntryMemA_line_words_1_MPORT_en & cacheEntryMemA_line_words_1_MPORT_mask) begin
      cacheEntryMemA_line_words_1[cacheEntryMemA_line_words_1_MPORT_addr] <= cacheEntryMemA_line_words_1_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[8:2];
    end
    if (cacheEntryMemA_line_words_2_MPORT_en & cacheEntryMemA_line_words_2_MPORT_mask) begin
      cacheEntryMemA_line_words_2[cacheEntryMemA_line_words_2_MPORT_addr] <= cacheEntryMemA_line_words_2_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[8:2];
    end
    if (cacheEntryMemA_line_words_3_MPORT_en & cacheEntryMemA_line_words_3_MPORT_mask) begin
      cacheEntryMemA_line_words_3[cacheEntryMemA_line_words_3_MPORT_addr] <= cacheEntryMemA_line_words_3_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[8:2];
    end
    if (cacheEntryMemB_valid_MPORT_1_en & cacheEntryMemB_valid_MPORT_1_mask) begin
      cacheEntryMemB_valid[cacheEntryMemB_valid_MPORT_1_addr] <= cacheEntryMemB_valid_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_valid_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_valid_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[8:2];
    end
    if (cacheEntryMemB_tag_MPORT_1_en & cacheEntryMemB_tag_MPORT_1_mask) begin
      cacheEntryMemB_tag[cacheEntryMemB_tag_MPORT_1_addr] <= cacheEntryMemB_tag_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_tag_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_tag_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[8:2];
    end
    if (cacheEntryMemB_line_words_0_MPORT_1_en & cacheEntryMemB_line_words_0_MPORT_1_mask) begin
      cacheEntryMemB_line_words_0[cacheEntryMemB_line_words_0_MPORT_1_addr] <= cacheEntryMemB_line_words_0_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[8:2];
    end
    if (cacheEntryMemB_line_words_1_MPORT_1_en & cacheEntryMemB_line_words_1_MPORT_1_mask) begin
      cacheEntryMemB_line_words_1[cacheEntryMemB_line_words_1_MPORT_1_addr] <= cacheEntryMemB_line_words_1_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[8:2];
    end
    if (cacheEntryMemB_line_words_2_MPORT_1_en & cacheEntryMemB_line_words_2_MPORT_1_mask) begin
      cacheEntryMemB_line_words_2[cacheEntryMemB_line_words_2_MPORT_1_addr] <= cacheEntryMemB_line_words_2_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[8:2];
    end
    if (cacheEntryMemB_line_words_3_MPORT_1_en & cacheEntryMemB_line_words_3_MPORT_1_mask) begin
      cacheEntryMemB_line_words_3[cacheEntryMemB_line_words_3_MPORT_1_addr] <= cacheEntryMemB_line_words_3_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[8:2];
    end
    if (reset) begin // @[ReadCache.scala 84:25]
      stateReg <= 3'h0; // @[ReadCache.scala 84:25]
    end else if (3'h0 == stateReg) begin // @[ReadCache.scala 194:20]
      if (initCounterWrap) begin // @[ReadCache.scala 197:29]
        stateReg <= 3'h1; // @[ReadCache.scala 197:40]
      end
    end else if (3'h1 == stateReg) begin // @[ReadCache.scala 194:20]
      if (start) begin // @[ReadCache.scala 202:19]
        stateReg <= 3'h2; // @[ReadCache.scala 202:30]
      end
    end else if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
      stateReg <= _GEN_72;
    end else begin
      stateReg <= _GEN_81;
    end
    if (start) begin // @[Reg.scala 20:18]
      offsetReg <= offsetReg_offset; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_rd <= io_in_rd; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_addr_tag <= request_addr_tag; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_addr_index <= request_addr_index; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_addr_offset <= request_addr_offset; // @[Reg.scala 20:22]
    end
    if (3'h0 == stateReg) begin // @[ReadCache.scala 194:20]
      doutReg <= _GEN_58;
    end else if (3'h1 == stateReg) begin // @[ReadCache.scala 194:20]
      doutReg <= _GEN_58;
    end else if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
      if (hit) begin // @[ReadCache.scala 207:17]
        doutReg <= _doutReg_T_9; // @[ReadCache.scala 182:13]
      end else begin
        doutReg <= _GEN_58;
      end
    end else begin
      doutReg <= _GEN_58;
    end
    if (3'h0 == stateReg) begin // @[ReadCache.scala 194:20]
      validReg <= _GEN_59;
    end else if (3'h1 == stateReg) begin // @[ReadCache.scala 194:20]
      validReg <= _GEN_59;
    end else if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
      validReg <= _GEN_74;
    end else begin
      validReg <= _GEN_59;
    end
    if (!(3'h0 == stateReg)) begin // @[ReadCache.scala 194:20]
      if (!(3'h1 == stateReg)) begin // @[ReadCache.scala 194:20]
        if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
          if (hit) begin // @[ReadCache.scala 207:17]
            lruReg <= _lruReg_T_5; // @[ReadCache.scala 184:12]
          end else begin
            lruReg <= _GEN_71;
          end
        end
      end
    end
    if (3'h0 == stateReg) begin // @[ReadCache.scala 194:20]
      wayReg <= _nextWay_T_2; // @[ReadCache.scala 169:11]
    end else if (3'h1 == stateReg) begin // @[ReadCache.scala 194:20]
      wayReg <= _nextWay_T_2; // @[ReadCache.scala 169:11]
    end else if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
      if (hit) begin // @[ReadCache.scala 207:17]
        wayReg <= ~hitA; // @[ReadCache.scala 185:13]
      end else begin
        wayReg <= _nextWay_T_2; // @[ReadCache.scala 169:11]
      end
    end else begin
      wayReg <= _nextWay_T_2; // @[ReadCache.scala 169:11]
    end
    cacheEntryReg_valid <= burstCounterEnable | _GEN_10; // @[ReadCache.scala 172:53 175:19]
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      cacheEntryReg_tag <= requestReg_addr_tag; // @[ReadCache.scala 175:19]
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_tag <= cacheEntryMemB_tag_cacheEntryB_data;
      end else begin
        cacheEntryReg_tag <= cacheEntryMemA_tag_cacheEntryA_data;
      end
    end
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      if (2'h0 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_0 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_line_words_0 <= cacheEntryMemB_line_words_0_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_0 <= cacheEntryMemA_line_words_0_cacheEntryA_data;
      end
    end
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      if (2'h1 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_1 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_line_words_1 <= cacheEntryMemB_line_words_1_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_1 <= cacheEntryMemA_line_words_1_cacheEntryA_data;
      end
    end
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      if (2'h2 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_2 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_line_words_2 <= cacheEntryMemB_line_words_2_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_2 <= cacheEntryMemA_line_words_2_cacheEntryA_data;
      end
    end
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      if (2'h3 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_3 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_line_words_3 <= cacheEntryMemB_line_words_3_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_3 <= cacheEntryMemA_line_words_3_cacheEntryA_data;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      initCounter <= 7'h0; // @[Counter.scala 61:40]
    end else if (_T) begin // @[Counter.scala 118:16]
      initCounter <= _wrap_value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      burstCounter <= 2'h0; // @[Counter.scala 61:40]
    end else if (burstCounterEnable) begin // @[Counter.scala 118:16]
      burstCounter <= _wrap_value_T_3; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cacheEntryMemA_valid[initvar] = _RAND_0[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cacheEntryMemA_tag[initvar] = _RAND_3[10:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cacheEntryMemA_line_words_0[initvar] = _RAND_6[15:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cacheEntryMemA_line_words_1[initvar] = _RAND_9[15:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cacheEntryMemA_line_words_2[initvar] = _RAND_12[15:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cacheEntryMemA_line_words_3[initvar] = _RAND_15[15:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cacheEntryMemB_valid[initvar] = _RAND_18[0:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cacheEntryMemB_tag[initvar] = _RAND_21[10:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cacheEntryMemB_line_words_0[initvar] = _RAND_24[15:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cacheEntryMemB_line_words_1[initvar] = _RAND_27[15:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cacheEntryMemB_line_words_2[initvar] = _RAND_30[15:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cacheEntryMemB_line_words_3[initvar] = _RAND_33[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cacheEntryMemA_valid_cacheEntryA_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cacheEntryMemA_valid_cacheEntryA_addr_pipe_0 = _RAND_2[6:0];
  _RAND_4 = {1{`RANDOM}};
  cacheEntryMemA_tag_cacheEntryA_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cacheEntryMemA_tag_cacheEntryA_addr_pipe_0 = _RAND_5[6:0];
  _RAND_7 = {1{`RANDOM}};
  cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0 = _RAND_8[6:0];
  _RAND_10 = {1{`RANDOM}};
  cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0 = _RAND_11[6:0];
  _RAND_13 = {1{`RANDOM}};
  cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0 = _RAND_14[6:0];
  _RAND_16 = {1{`RANDOM}};
  cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0 = _RAND_17[6:0];
  _RAND_19 = {1{`RANDOM}};
  cacheEntryMemB_valid_cacheEntryB_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  cacheEntryMemB_valid_cacheEntryB_addr_pipe_0 = _RAND_20[6:0];
  _RAND_22 = {1{`RANDOM}};
  cacheEntryMemB_tag_cacheEntryB_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  cacheEntryMemB_tag_cacheEntryB_addr_pipe_0 = _RAND_23[6:0];
  _RAND_25 = {1{`RANDOM}};
  cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0 = _RAND_26[6:0];
  _RAND_28 = {1{`RANDOM}};
  cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0 = _RAND_29[6:0];
  _RAND_31 = {1{`RANDOM}};
  cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0 = _RAND_32[6:0];
  _RAND_34 = {1{`RANDOM}};
  cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0 = _RAND_35[6:0];
  _RAND_36 = {1{`RANDOM}};
  stateReg = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  offsetReg = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  requestReg_rd = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  requestReg_addr_tag = _RAND_39[10:0];
  _RAND_40 = {1{`RANDOM}};
  requestReg_addr_index = _RAND_40[6:0];
  _RAND_41 = {1{`RANDOM}};
  requestReg_addr_offset = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  doutReg = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  validReg = _RAND_43[0:0];
  _RAND_44 = {4{`RANDOM}};
  lruReg = _RAND_44[127:0];
  _RAND_45 = {1{`RANDOM}};
  wayReg = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  cacheEntryReg_valid = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  cacheEntryReg_tag = _RAND_47[10:0];
  _RAND_48 = {1{`RANDOM}};
  cacheEntryReg_line_words_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  cacheEntryReg_line_words_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  cacheEntryReg_line_words_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  cacheEntryReg_line_words_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  initCounter = _RAND_52[6:0];
  _RAND_53 = {1{`RANDOM}};
  burstCounter = _RAND_53[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cache(
  input         clock,
  input         reset,
  input         io_enable,
  input         io_in_rd,
  input         io_in_wr,
  input  [6:0]  io_in_addr,
  input  [15:0] io_in_din,
  output [15:0] io_in_dout,
  output        io_in_wait_n,
  output        io_in_valid,
  output        io_out_rd,
  output        io_out_wr,
  output [24:0] io_out_addr,
  output [15:0] io_out_din,
  input  [15:0] io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_39;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
`endif // RANDOMIZE_REG_INIT
  reg  cacheEntryMemA_valid [0:1]; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_valid_cacheEntryA_en; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_valid_cacheEntryA_addr; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_valid_cacheEntryA_data; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_valid_MPORT_data; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_valid_MPORT_addr; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_valid_MPORT_mask; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_valid_MPORT_en; // @[Cache.scala 115:35]
  reg  cacheEntryMemA_valid_cacheEntryA_en_pipe_0;
  reg  cacheEntryMemA_valid_cacheEntryA_addr_pipe_0;
  reg  cacheEntryMemA_dirty [0:1]; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_dirty_cacheEntryA_en; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_dirty_cacheEntryA_addr; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_dirty_cacheEntryA_data; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_dirty_MPORT_data; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_dirty_MPORT_addr; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_dirty_MPORT_mask; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_dirty_MPORT_en; // @[Cache.scala 115:35]
  reg  cacheEntryMemA_dirty_cacheEntryA_en_pipe_0;
  reg  cacheEntryMemA_dirty_cacheEntryA_addr_pipe_0;
  reg [3:0] cacheEntryMemA_tag [0:1]; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_tag_cacheEntryA_en; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_tag_cacheEntryA_addr; // @[Cache.scala 115:35]
  wire [3:0] cacheEntryMemA_tag_cacheEntryA_data; // @[Cache.scala 115:35]
  wire [3:0] cacheEntryMemA_tag_MPORT_data; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_tag_MPORT_addr; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_tag_MPORT_mask; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_tag_MPORT_en; // @[Cache.scala 115:35]
  reg  cacheEntryMemA_tag_cacheEntryA_en_pipe_0;
  reg  cacheEntryMemA_tag_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_0 [0:1]; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_0_cacheEntryA_en; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_0_cacheEntryA_addr; // @[Cache.scala 115:35]
  wire [15:0] cacheEntryMemA_line_words_0_cacheEntryA_data; // @[Cache.scala 115:35]
  wire [15:0] cacheEntryMemA_line_words_0_MPORT_data; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_0_MPORT_addr; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_0_MPORT_mask; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_0_MPORT_en; // @[Cache.scala 115:35]
  reg  cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0;
  reg  cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_1 [0:1]; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_1_cacheEntryA_en; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_1_cacheEntryA_addr; // @[Cache.scala 115:35]
  wire [15:0] cacheEntryMemA_line_words_1_cacheEntryA_data; // @[Cache.scala 115:35]
  wire [15:0] cacheEntryMemA_line_words_1_MPORT_data; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_1_MPORT_addr; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_1_MPORT_mask; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_1_MPORT_en; // @[Cache.scala 115:35]
  reg  cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0;
  reg  cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_2 [0:1]; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_2_cacheEntryA_en; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_2_cacheEntryA_addr; // @[Cache.scala 115:35]
  wire [15:0] cacheEntryMemA_line_words_2_cacheEntryA_data; // @[Cache.scala 115:35]
  wire [15:0] cacheEntryMemA_line_words_2_MPORT_data; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_2_MPORT_addr; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_2_MPORT_mask; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_2_MPORT_en; // @[Cache.scala 115:35]
  reg  cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0;
  reg  cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_3 [0:1]; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_3_cacheEntryA_en; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_3_cacheEntryA_addr; // @[Cache.scala 115:35]
  wire [15:0] cacheEntryMemA_line_words_3_cacheEntryA_data; // @[Cache.scala 115:35]
  wire [15:0] cacheEntryMemA_line_words_3_MPORT_data; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_3_MPORT_addr; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_3_MPORT_mask; // @[Cache.scala 115:35]
  wire  cacheEntryMemA_line_words_3_MPORT_en; // @[Cache.scala 115:35]
  reg  cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0;
  reg  cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0;
  reg  cacheEntryMemB_valid [0:1]; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_valid_cacheEntryB_en; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_valid_cacheEntryB_addr; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_valid_cacheEntryB_data; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_valid_MPORT_1_data; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_valid_MPORT_1_addr; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_valid_MPORT_1_mask; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_valid_MPORT_1_en; // @[Cache.scala 116:35]
  reg  cacheEntryMemB_valid_cacheEntryB_en_pipe_0;
  reg  cacheEntryMemB_valid_cacheEntryB_addr_pipe_0;
  reg  cacheEntryMemB_dirty [0:1]; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_dirty_cacheEntryB_en; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_dirty_cacheEntryB_addr; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_dirty_cacheEntryB_data; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_dirty_MPORT_1_data; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_dirty_MPORT_1_addr; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_dirty_MPORT_1_mask; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_dirty_MPORT_1_en; // @[Cache.scala 116:35]
  reg  cacheEntryMemB_dirty_cacheEntryB_en_pipe_0;
  reg  cacheEntryMemB_dirty_cacheEntryB_addr_pipe_0;
  reg [3:0] cacheEntryMemB_tag [0:1]; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_tag_cacheEntryB_en; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_tag_cacheEntryB_addr; // @[Cache.scala 116:35]
  wire [3:0] cacheEntryMemB_tag_cacheEntryB_data; // @[Cache.scala 116:35]
  wire [3:0] cacheEntryMemB_tag_MPORT_1_data; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_tag_MPORT_1_addr; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_tag_MPORT_1_mask; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_tag_MPORT_1_en; // @[Cache.scala 116:35]
  reg  cacheEntryMemB_tag_cacheEntryB_en_pipe_0;
  reg  cacheEntryMemB_tag_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_0 [0:1]; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_0_cacheEntryB_en; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_0_cacheEntryB_addr; // @[Cache.scala 116:35]
  wire [15:0] cacheEntryMemB_line_words_0_cacheEntryB_data; // @[Cache.scala 116:35]
  wire [15:0] cacheEntryMemB_line_words_0_MPORT_1_data; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_0_MPORT_1_addr; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_0_MPORT_1_mask; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_0_MPORT_1_en; // @[Cache.scala 116:35]
  reg  cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0;
  reg  cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_1 [0:1]; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_1_cacheEntryB_en; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_1_cacheEntryB_addr; // @[Cache.scala 116:35]
  wire [15:0] cacheEntryMemB_line_words_1_cacheEntryB_data; // @[Cache.scala 116:35]
  wire [15:0] cacheEntryMemB_line_words_1_MPORT_1_data; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_1_MPORT_1_addr; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_1_MPORT_1_mask; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_1_MPORT_1_en; // @[Cache.scala 116:35]
  reg  cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0;
  reg  cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_2 [0:1]; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_2_cacheEntryB_en; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_2_cacheEntryB_addr; // @[Cache.scala 116:35]
  wire [15:0] cacheEntryMemB_line_words_2_cacheEntryB_data; // @[Cache.scala 116:35]
  wire [15:0] cacheEntryMemB_line_words_2_MPORT_1_data; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_2_MPORT_1_addr; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_2_MPORT_1_mask; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_2_MPORT_1_en; // @[Cache.scala 116:35]
  reg  cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0;
  reg  cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_3 [0:1]; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_3_cacheEntryB_en; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_3_cacheEntryB_addr; // @[Cache.scala 116:35]
  wire [15:0] cacheEntryMemB_line_words_3_cacheEntryB_data; // @[Cache.scala 116:35]
  wire [15:0] cacheEntryMemB_line_words_3_MPORT_1_data; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_3_MPORT_1_addr; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_3_MPORT_1_mask; // @[Cache.scala 116:35]
  wire  cacheEntryMemB_line_words_3_MPORT_1_en; // @[Cache.scala 116:35]
  reg  cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0;
  reg  cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0;
  reg [3:0] stateReg; // @[Cache.scala 87:25]
  wire [5:0] offsetReg_addr = io_in_addr[6:1]; // @[Cache.scala 94:27]
  wire [1:0] offsetReg_offset = offsetReg_addr[1:0]; // @[Cache.scala 95:22]
  reg [1:0] offsetReg; // @[Reg.scala 19:16]
  wire  _start_T_2 = stateReg == 4'h1; // @[Cache.scala 149:64]
  wire  start = io_enable & (io_in_rd | io_in_wr) & stateReg == 4'h1; // @[Cache.scala 149:52]
  wire [6:0] _request_WIRE_1 = {{1'd0}, offsetReg_addr};
  wire [1:0] request_addr_offset = _request_WIRE_1[1:0]; // @[Address.scala 78:49]
  wire  request_addr_index = _request_WIRE_1[2]; // @[Address.scala 78:49]
  wire [3:0] request_addr_tag = _request_WIRE_1[6:3]; // @[Address.scala 78:49]
  reg  requestReg_rd; // @[Reg.scala 19:16]
  reg  requestReg_wr; // @[Reg.scala 19:16]
  reg [3:0] requestReg_addr_tag; // @[Reg.scala 19:16]
  reg  requestReg_addr_index; // @[Reg.scala 19:16]
  reg [1:0] requestReg_addr_offset; // @[Reg.scala 19:16]
  reg [15:0] requestReg_din; // @[Reg.scala 19:16]
  reg [15:0] doutReg; // @[Cache.scala 104:20]
  reg  validReg; // @[Cache.scala 105:25]
  reg [1:0] lruReg; // @[Cache.scala 108:19]
  reg  wayReg; // @[Cache.scala 112:23]
  wire [1:0] _nextWay_T = lruReg >> request_addr_index; // @[Cache.scala 181:31]
  wire  _nextWay_T_2 = start ? _nextWay_T[0] : wayReg; // @[Cache.scala 181:17]
  wire  hitA = cacheEntryMemA_valid_cacheEntryA_data & cacheEntryMemA_tag_cacheEntryA_data == requestReg_addr_tag; // @[Entry.scala 59:42]
  wire  hitB = cacheEntryMemB_valid_cacheEntryB_data & cacheEntryMemB_tag_cacheEntryB_data == requestReg_addr_tag; // @[Entry.scala 59:42]
  wire  hit = hitA | hitB; // @[Cache.scala 153:18]
  wire  _GEN_96 = hit ? ~hitA : _nextWay_T_2; // @[Cache.scala 181:11 207:13 234:17]
  wire  _GEN_111 = 4'h2 == stateReg ? _GEN_96 : _nextWay_T_2; // @[Cache.scala 181:11 221:20]
  wire  _GEN_116 = 4'h1 == stateReg ? _nextWay_T_2 : _GEN_111; // @[Cache.scala 181:11 221:20]
  wire  nextWay = 4'h0 == stateReg ? _nextWay_T_2 : _GEN_116; // @[Cache.scala 181:11 221:20]
  wire  _cacheEntryReg_T_valid = nextWay ? cacheEntryMemB_valid_cacheEntryB_data : cacheEntryMemA_valid_cacheEntryA_data
    ; // @[Cache.scala 124:36]
  wire  _cacheEntryReg_T_dirty = nextWay ? cacheEntryMemB_dirty_cacheEntryB_data : cacheEntryMemA_dirty_cacheEntryA_data
    ; // @[Cache.scala 124:36]
  wire  _cacheEntryReg_T_1 = stateReg == 4'h2; // @[Cache.scala 124:82]
  reg  cacheEntryReg_valid; // @[Reg.scala 19:16]
  reg  cacheEntryReg_dirty; // @[Reg.scala 19:16]
  reg [3:0] cacheEntryReg_tag; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_0; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_1; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_2; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_3; // @[Reg.scala 19:16]
  wire  _GEN_13 = _cacheEntryReg_T_1 ? _cacheEntryReg_T_valid : cacheEntryReg_valid; // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_14 = _cacheEntryReg_T_1 ? _cacheEntryReg_T_dirty : cacheEntryReg_dirty; // @[Reg.scala 19:16 20:{18,22}]
  wire  _nextCacheEntry_T = stateReg == 4'h8; // @[Cache.scala 127:37]
  wire  _T = stateReg == 4'h0; // @[Cache.scala 129:17]
  wire  _T_2 = ~wayReg; // @[Cache.scala 129:64]
  wire  _T_3 = _nextCacheEntry_T & ~wayReg; // @[Cache.scala 129:61]
  wire  _T_7 = _nextCacheEntry_T & wayReg; // @[Cache.scala 133:61]
  wire  burstCounterEnable_fill = stateReg == 4'h4 & io_out_valid; // @[Cache.scala 139:44]
  wire  _burstCounterEnable_evict_T = stateReg == 4'h5; // @[Cache.scala 140:27]
  wire  _burstCounterEnable_evict_T_1 = stateReg == 4'h6; // @[Cache.scala 140:55]
  wire  burstCounterEnable_evict = (stateReg == 4'h5 | stateReg == 4'h6) & io_out_wait_n; // @[Cache.scala 140:76]
  wire  burstCounterEnable = burstCounterEnable_fill | burstCounterEnable_evict; // @[Cache.scala 141:10]
  reg  initCounter; // @[Counter.scala 61:40]
  wire  initCounterWrap = _T & initCounter; // @[Counter.scala 118:{16,23}]
  reg [1:0] burstCounter; // @[Counter.scala 61:40]
  wire  wrap_wrap_1 = burstCounter == 2'h3; // @[Counter.scala 73:24]
  wire [1:0] _wrap_value_T_3 = burstCounter + 2'h1; // @[Counter.scala 77:24]
  wire  burstCounterWrap = burstCounterEnable & wrap_wrap_1; // @[Counter.scala 118:{16,23}]
  wire  miss = ~hit; // @[Cache.scala 154:14]
  wire  dirtyA = cacheEntryMemA_dirty_cacheEntryA_data & cacheEntryMemA_tag_cacheEntryA_data != requestReg_addr_tag; // @[Entry.scala 66:44]
  wire  dirtyB = cacheEntryMemB_dirty_cacheEntryB_data & cacheEntryMemB_tag_cacheEntryB_data != requestReg_addr_tag; // @[Entry.scala 66:44]
  wire  dirty = _T_2 & dirtyA | wayReg & dirtyB; // @[Cache.scala 157:35]
  wire  wordDone = burstCounter == 2'h0; // @[Cache.scala 163:18]
  wire [3:0] _outAddr_addr_T_1_tag = stateReg == 4'h3 ? requestReg_addr_tag : cacheEntryReg_tag; // @[Cache.scala 176:19]
  wire [1:0] _outAddr_addr_T_1_offset = stateReg == 4'h3 ? requestReg_addr_offset : 2'h0; // @[Cache.scala 176:19]
  wire [6:0] outAddr_addr = {_outAddr_addr_T_1_tag,requestReg_addr_index,_outAddr_addr_T_1_offset}; // @[Cache.scala 176:66]
  wire [7:0] outAddr = {outAddr_addr, 1'h0}; // @[Cache.scala 177:11]
  wire [1:0] n = requestReg_addr_offset + burstCounter; // @[Cache.scala 185:57]
  wire [15:0] entry_line_words_0 = 2'h0 == n ? io_out_dout : cacheEntryReg_line_words_0; // @[Entry.scala 92:11 93:{30,30}]
  wire [15:0] entry_line_words_1 = 2'h1 == n ? io_out_dout : cacheEntryReg_line_words_1; // @[Entry.scala 92:11 93:{30,30}]
  wire [15:0] entry_line_words_2 = 2'h2 == n ? io_out_dout : cacheEntryReg_line_words_2; // @[Entry.scala 92:11 93:{30,30}]
  wire [15:0] entry_line_words_3 = 2'h3 == n ? io_out_dout : cacheEntryReg_line_words_3; // @[Entry.scala 92:11 93:{30,30}]
  wire [63:0] _doutReg_ws_T = {entry_line_words_3,entry_line_words_2,entry_line_words_1,entry_line_words_0}; // @[Line.scala 77:32]
  wire [15:0] doutReg_ws_0 = _doutReg_ws_T[15:0]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_1 = _doutReg_ws_T[31:16]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_2 = _doutReg_ws_T[47:32]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_3 = _doutReg_ws_T[63:48]; // @[Util.scala 104:11]
  wire [15:0] _GEN_51 = 2'h1 == offsetReg ? doutReg_ws_1 : doutReg_ws_0; // @[Util.scala 104:{11,11}]
  wire [15:0] _GEN_52 = 2'h2 == offsetReg ? doutReg_ws_2 : _GEN_51; // @[Util.scala 104:{11,11}]
  wire [15:0] _GEN_53 = 2'h3 == offsetReg ? doutReg_ws_3 : _GEN_52; // @[Util.scala 104:{11,11}]
  wire [15:0] _doutReg_T_2 = {_GEN_53[7:0],_GEN_53[15:8]}; // @[Util.scala 114:49]
  wire  _GEN_54 = burstCounterEnable_fill | _GEN_13; // @[Cache.scala 184:53 187:19]
  wire  _GEN_55 = burstCounterEnable_fill ? cacheEntryReg_dirty : _GEN_14; // @[Cache.scala 184:53 187:19]
  wire [15:0] _GEN_61 = burstCounterEnable_fill ? _doutReg_T_2 : doutReg; // @[Cache.scala 184:53 188:13 104:20]
  wire  _GEN_62 = burstCounterEnable_fill & (requestReg_rd & wordDone); // @[Cache.scala 184:53 189:14 105:25]
  wire [63:0] _cacheEntryReg_words_ws_T = {cacheEntryReg_line_words_3,cacheEntryReg_line_words_2,
    cacheEntryReg_line_words_1,cacheEntryReg_line_words_0}; // @[Line.scala 77:32]
  wire [15:0] cacheEntryReg_words_ws_0 = _cacheEntryReg_words_ws_T[15:0]; // @[Util.scala 104:11]
  wire [15:0] cacheEntryReg_words_ws_1 = _cacheEntryReg_words_ws_T[31:16]; // @[Util.scala 104:11]
  wire [15:0] cacheEntryReg_words_ws_2 = _cacheEntryReg_words_ws_T[47:32]; // @[Util.scala 104:11]
  wire [15:0] cacheEntryReg_words_ws_3 = _cacheEntryReg_words_ws_T[63:48]; // @[Util.scala 104:11]
  wire [15:0] _cacheEntryReg_words_T_2 = {requestReg_din[7:0],requestReg_din[15:8]}; // @[Util.scala 114:49]
  wire [15:0] cacheEntryReg_words_0 = 2'h0 == offsetReg ? _cacheEntryReg_words_T_2 : cacheEntryReg_words_ws_0; // @[Entry.scala 108:{19,19}]
  wire [15:0] cacheEntryReg_words_1 = 2'h1 == offsetReg ? _cacheEntryReg_words_T_2 : cacheEntryReg_words_ws_1; // @[Entry.scala 108:{19,19}]
  wire [15:0] cacheEntryReg_words_2 = 2'h2 == offsetReg ? _cacheEntryReg_words_T_2 : cacheEntryReg_words_ws_2; // @[Entry.scala 108:{19,19}]
  wire [15:0] cacheEntryReg_words_3 = 2'h3 == offsetReg ? _cacheEntryReg_words_T_2 : cacheEntryReg_words_ws_3; // @[Entry.scala 108:{19,19}]
  wire [63:0] _cacheEntryReg_T_2 = {cacheEntryReg_words_3,cacheEntryReg_words_2,cacheEntryReg_words_1,
    cacheEntryReg_words_0}; // @[Entry.scala 112:39]
  wire [15:0] cacheEntryReg_entry_line_words_0 = _cacheEntryReg_T_2[15:0]; // @[Entry.scala 112:39]
  wire [15:0] cacheEntryReg_entry_line_words_1 = _cacheEntryReg_T_2[31:16]; // @[Entry.scala 112:39]
  wire [15:0] cacheEntryReg_entry_line_words_2 = _cacheEntryReg_T_2[47:32]; // @[Entry.scala 112:39]
  wire [15:0] cacheEntryReg_entry_line_words_3 = _cacheEntryReg_T_2[63:48]; // @[Entry.scala 112:39]
  wire [3:0] _GEN_67 = stateReg == 4'h7 ? 4'h8 : stateReg; // @[Cache.scala 193:34 194:14 87:25]
  wire [63:0] _doutReg_ws_T_1 = {cacheEntryMemA_line_words_3_cacheEntryA_data,
    cacheEntryMemA_line_words_2_cacheEntryA_data,cacheEntryMemA_line_words_1_cacheEntryA_data,
    cacheEntryMemA_line_words_0_cacheEntryA_data}; // @[Line.scala 77:32]
  wire [15:0] doutReg_ws_0_1 = _doutReg_ws_T_1[15:0]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_1_1 = _doutReg_ws_T_1[31:16]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_2_1 = _doutReg_ws_T_1[47:32]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_3_1 = _doutReg_ws_T_1[63:48]; // @[Util.scala 104:11]
  wire [15:0] _GEN_78 = 2'h1 == offsetReg ? doutReg_ws_1_1 : doutReg_ws_0_1; // @[Util.scala 104:{11,11}]
  wire [15:0] _GEN_79 = 2'h2 == offsetReg ? doutReg_ws_2_1 : _GEN_78; // @[Util.scala 104:{11,11}]
  wire [15:0] _GEN_80 = 2'h3 == offsetReg ? doutReg_ws_3_1 : _GEN_79; // @[Util.scala 104:{11,11}]
  wire [15:0] _doutReg_T_5 = {_GEN_80[7:0],_GEN_80[15:8]}; // @[Util.scala 114:49]
  wire [63:0] _doutReg_ws_T_2 = {cacheEntryMemB_line_words_3_cacheEntryB_data,
    cacheEntryMemB_line_words_2_cacheEntryB_data,cacheEntryMemB_line_words_1_cacheEntryB_data,
    cacheEntryMemB_line_words_0_cacheEntryB_data}; // @[Line.scala 77:32]
  wire [15:0] doutReg_ws_0_2 = _doutReg_ws_T_2[15:0]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_1_2 = _doutReg_ws_T_2[31:16]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_2_2 = _doutReg_ws_T_2[47:32]; // @[Util.scala 104:11]
  wire [15:0] doutReg_ws_3_2 = _doutReg_ws_T_2[63:48]; // @[Util.scala 104:11]
  wire [15:0] _GEN_82 = 2'h1 == offsetReg ? doutReg_ws_1_2 : doutReg_ws_0_2; // @[Util.scala 104:{11,11}]
  wire [15:0] _GEN_83 = 2'h2 == offsetReg ? doutReg_ws_2_2 : _GEN_82; // @[Util.scala 104:{11,11}]
  wire [15:0] _GEN_84 = 2'h3 == offsetReg ? doutReg_ws_3_2 : _GEN_83; // @[Util.scala 104:{11,11}]
  wire [15:0] _doutReg_T_8 = {_GEN_84[7:0],_GEN_84[15:8]}; // @[Util.scala 114:49]
  wire [15:0] _doutReg_T_9 = hitA ? _doutReg_T_5 : _doutReg_T_8; // @[Cache.scala 201:21]
  wire [3:0] _GEN_85 = requestReg_rd ? 4'h1 : 4'h7; // @[Cache.scala 199:25 200:16 204:16]
  wire [15:0] _GEN_86 = requestReg_rd ? _doutReg_T_9 : _GEN_61; // @[Cache.scala 199:25 201:15]
  wire  _GEN_87 = requestReg_rd | _GEN_62; // @[Cache.scala 199:25 202:16]
  wire [1:0] _lruReg_T = 2'h1 << requestReg_addr_index; // @[Cache.scala 206:28]
  wire [1:0] _lruReg_T_1 = lruReg | _lruReg_T; // @[Cache.scala 206:28]
  wire [1:0] _lruReg_T_2 = ~lruReg; // @[Cache.scala 206:28]
  wire [1:0] _lruReg_T_3 = _lruReg_T_2 | _lruReg_T; // @[Cache.scala 206:28]
  wire [1:0] _lruReg_T_4 = ~_lruReg_T_3; // @[Cache.scala 206:28]
  wire [1:0] _lruReg_T_5 = hitA ? _lruReg_T_1 : _lruReg_T_4; // @[Cache.scala 206:28]
  wire [1:0] _lruReg_T_12 = _T_2 ? _lruReg_T_1 : _lruReg_T_4; // @[Cache.scala 217:28]
  wire [3:0] _GEN_88 = miss ? 4'h3 : _GEN_67; // @[Cache.scala 211:14 234:74]
  wire [1:0] _GEN_89 = miss ? _lruReg_T_12 : lruReg; // @[Cache.scala 212:12 108:19 234:74]
  wire [3:0] _GEN_90 = dirty ? 4'h5 : _GEN_88; // @[Cache.scala 216:14 234:45]
  wire [1:0] _GEN_91 = dirty ? _lruReg_T_12 : _GEN_89; // @[Cache.scala 217:12 234:45]
  wire [3:0] _GEN_92 = hit ? _GEN_85 : _GEN_90; // @[Cache.scala 234:17]
  wire [3:0] _GEN_97 = io_out_wait_n ? 4'h4 : _GEN_67; // @[Cache.scala 239:{27,38}]
  wire [3:0] _stateReg_T = requestReg_wr ? 4'h7 : 4'h8; // @[Cache.scala 245:24]
  wire [3:0] _GEN_98 = burstCounterWrap ? _stateReg_T : _GEN_67; // @[Cache.scala 244:30 245:18]
  wire [3:0] _GEN_99 = io_out_wait_n ? 4'h6 : _GEN_67; // @[Cache.scala 251:{27,38}]
  wire [3:0] _GEN_100 = burstCounterWrap ? 4'h3 : _GEN_67; // @[Cache.scala 256:{30,41}]
  wire [3:0] _GEN_101 = 4'h8 == stateReg ? 4'h1 : _GEN_67; // @[Cache.scala 221:20 263:32]
  wire [3:0] _GEN_102 = 4'h7 == stateReg ? 4'h8 : _GEN_101; // @[Cache.scala 221:20 260:32]
  wire [3:0] _GEN_103 = 4'h6 == stateReg ? _GEN_100 : _GEN_102; // @[Cache.scala 221:20]
  wire [3:0] _GEN_104 = 4'h5 == stateReg ? _GEN_99 : _GEN_103; // @[Cache.scala 221:20]
  wire [3:0] _GEN_105 = 4'h4 == stateReg ? _GEN_98 : _GEN_104; // @[Cache.scala 221:20]
  wire [3:0] _GEN_106 = 4'h3 == stateReg ? _GEN_97 : _GEN_105; // @[Cache.scala 221:20]
  wire [15:0] _GEN_123 = 2'h1 == burstCounter ? cacheEntryReg_line_words_1 : cacheEntryReg_line_words_0; // @[Cache.scala 275:{14,14}]
  wire [15:0] _GEN_124 = 2'h2 == burstCounter ? cacheEntryReg_line_words_2 : _GEN_123; // @[Cache.scala 275:{14,14}]
  assign cacheEntryMemA_valid_cacheEntryA_en = cacheEntryMemA_valid_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_valid_cacheEntryA_addr = cacheEntryMemA_valid_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_valid_cacheEntryA_data = cacheEntryMemA_valid[cacheEntryMemA_valid_cacheEntryA_addr]; // @[Cache.scala 115:35]
  assign cacheEntryMemA_valid_MPORT_data = _nextCacheEntry_T & cacheEntryReg_valid;
  assign cacheEntryMemA_valid_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_valid_MPORT_mask = 1'h1;
  assign cacheEntryMemA_valid_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_dirty_cacheEntryA_en = cacheEntryMemA_dirty_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_dirty_cacheEntryA_addr = cacheEntryMemA_dirty_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_dirty_cacheEntryA_data = cacheEntryMemA_dirty[cacheEntryMemA_dirty_cacheEntryA_addr]; // @[Cache.scala 115:35]
  assign cacheEntryMemA_dirty_MPORT_data = _nextCacheEntry_T & cacheEntryReg_dirty;
  assign cacheEntryMemA_dirty_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_dirty_MPORT_mask = 1'h1;
  assign cacheEntryMemA_dirty_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_tag_cacheEntryA_en = cacheEntryMemA_tag_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_tag_cacheEntryA_addr = cacheEntryMemA_tag_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_tag_cacheEntryA_data = cacheEntryMemA_tag[cacheEntryMemA_tag_cacheEntryA_addr]; // @[Cache.scala 115:35]
  assign cacheEntryMemA_tag_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_tag : 4'h0;
  assign cacheEntryMemA_tag_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_tag_MPORT_mask = 1'h1;
  assign cacheEntryMemA_tag_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_0_cacheEntryA_en = cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_0_cacheEntryA_addr = cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_0_cacheEntryA_data =
    cacheEntryMemA_line_words_0[cacheEntryMemA_line_words_0_cacheEntryA_addr]; // @[Cache.scala 115:35]
  assign cacheEntryMemA_line_words_0_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_0 : 16'h0;
  assign cacheEntryMemA_line_words_0_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_0_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_0_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_1_cacheEntryA_en = cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_1_cacheEntryA_addr = cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_1_cacheEntryA_data =
    cacheEntryMemA_line_words_1[cacheEntryMemA_line_words_1_cacheEntryA_addr]; // @[Cache.scala 115:35]
  assign cacheEntryMemA_line_words_1_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_1 : 16'h0;
  assign cacheEntryMemA_line_words_1_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_1_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_1_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_2_cacheEntryA_en = cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_2_cacheEntryA_addr = cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_2_cacheEntryA_data =
    cacheEntryMemA_line_words_2[cacheEntryMemA_line_words_2_cacheEntryA_addr]; // @[Cache.scala 115:35]
  assign cacheEntryMemA_line_words_2_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_2 : 16'h0;
  assign cacheEntryMemA_line_words_2_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_2_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_2_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_3_cacheEntryA_en = cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_3_cacheEntryA_addr = cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_3_cacheEntryA_data =
    cacheEntryMemA_line_words_3[cacheEntryMemA_line_words_3_cacheEntryA_addr]; // @[Cache.scala 115:35]
  assign cacheEntryMemA_line_words_3_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_3 : 16'h0;
  assign cacheEntryMemA_line_words_3_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_3_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_3_MPORT_en = _T | _T_3;
  assign cacheEntryMemB_valid_cacheEntryB_en = cacheEntryMemB_valid_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_valid_cacheEntryB_addr = cacheEntryMemB_valid_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_valid_cacheEntryB_data = cacheEntryMemB_valid[cacheEntryMemB_valid_cacheEntryB_addr]; // @[Cache.scala 116:35]
  assign cacheEntryMemB_valid_MPORT_1_data = _nextCacheEntry_T & cacheEntryReg_valid;
  assign cacheEntryMemB_valid_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_valid_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_valid_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_dirty_cacheEntryB_en = cacheEntryMemB_dirty_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_dirty_cacheEntryB_addr = cacheEntryMemB_dirty_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_dirty_cacheEntryB_data = cacheEntryMemB_dirty[cacheEntryMemB_dirty_cacheEntryB_addr]; // @[Cache.scala 116:35]
  assign cacheEntryMemB_dirty_MPORT_1_data = _nextCacheEntry_T & cacheEntryReg_dirty;
  assign cacheEntryMemB_dirty_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_dirty_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_dirty_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_tag_cacheEntryB_en = cacheEntryMemB_tag_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_tag_cacheEntryB_addr = cacheEntryMemB_tag_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_tag_cacheEntryB_data = cacheEntryMemB_tag[cacheEntryMemB_tag_cacheEntryB_addr]; // @[Cache.scala 116:35]
  assign cacheEntryMemB_tag_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_tag : 4'h0;
  assign cacheEntryMemB_tag_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_tag_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_tag_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_0_cacheEntryB_en = cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_0_cacheEntryB_addr = cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_0_cacheEntryB_data =
    cacheEntryMemB_line_words_0[cacheEntryMemB_line_words_0_cacheEntryB_addr]; // @[Cache.scala 116:35]
  assign cacheEntryMemB_line_words_0_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_0 : 16'h0;
  assign cacheEntryMemB_line_words_0_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_0_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_0_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_1_cacheEntryB_en = cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_1_cacheEntryB_addr = cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_1_cacheEntryB_data =
    cacheEntryMemB_line_words_1[cacheEntryMemB_line_words_1_cacheEntryB_addr]; // @[Cache.scala 116:35]
  assign cacheEntryMemB_line_words_1_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_1 : 16'h0;
  assign cacheEntryMemB_line_words_1_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_1_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_1_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_2_cacheEntryB_en = cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_2_cacheEntryB_addr = cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_2_cacheEntryB_data =
    cacheEntryMemB_line_words_2[cacheEntryMemB_line_words_2_cacheEntryB_addr]; // @[Cache.scala 116:35]
  assign cacheEntryMemB_line_words_2_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_2 : 16'h0;
  assign cacheEntryMemB_line_words_2_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_2_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_2_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_3_cacheEntryB_en = cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_3_cacheEntryB_addr = cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_3_cacheEntryB_data =
    cacheEntryMemB_line_words_3[cacheEntryMemB_line_words_3_cacheEntryB_addr]; // @[Cache.scala 116:35]
  assign cacheEntryMemB_line_words_3_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_3 : 16'h0;
  assign cacheEntryMemB_line_words_3_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_3_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_3_MPORT_1_en = _T | _T_7;
  assign io_in_dout = doutReg; // @[Cache.scala 269:14]
  assign io_in_wait_n = io_enable & _start_T_2; // @[Cache.scala 150:26]
  assign io_in_valid = validReg; // @[Cache.scala 268:15]
  assign io_out_rd = stateReg == 4'h3; // @[Cache.scala 270:25]
  assign io_out_wr = _burstCounterEnable_evict_T | _burstCounterEnable_evict_T_1; // @[Cache.scala 271:41]
  assign io_out_addr = {{17'd0}, outAddr}; // @[Cache.scala 273:15]
  assign io_out_din = 2'h3 == burstCounter ? cacheEntryReg_line_words_3 : _GEN_124; // @[Cache.scala 275:{14,14}]
  always @(posedge clock) begin
    if (cacheEntryMemA_valid_MPORT_en & cacheEntryMemA_valid_MPORT_mask) begin
      cacheEntryMemA_valid[cacheEntryMemA_valid_MPORT_addr] <= cacheEntryMemA_valid_MPORT_data; // @[Cache.scala 115:35]
    end
    cacheEntryMemA_valid_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_valid_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemA_dirty_MPORT_en & cacheEntryMemA_dirty_MPORT_mask) begin
      cacheEntryMemA_dirty[cacheEntryMemA_dirty_MPORT_addr] <= cacheEntryMemA_dirty_MPORT_data; // @[Cache.scala 115:35]
    end
    cacheEntryMemA_dirty_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_dirty_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemA_tag_MPORT_en & cacheEntryMemA_tag_MPORT_mask) begin
      cacheEntryMemA_tag[cacheEntryMemA_tag_MPORT_addr] <= cacheEntryMemA_tag_MPORT_data; // @[Cache.scala 115:35]
    end
    cacheEntryMemA_tag_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_tag_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemA_line_words_0_MPORT_en & cacheEntryMemA_line_words_0_MPORT_mask) begin
      cacheEntryMemA_line_words_0[cacheEntryMemA_line_words_0_MPORT_addr] <= cacheEntryMemA_line_words_0_MPORT_data; // @[Cache.scala 115:35]
    end
    cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemA_line_words_1_MPORT_en & cacheEntryMemA_line_words_1_MPORT_mask) begin
      cacheEntryMemA_line_words_1[cacheEntryMemA_line_words_1_MPORT_addr] <= cacheEntryMemA_line_words_1_MPORT_data; // @[Cache.scala 115:35]
    end
    cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemA_line_words_2_MPORT_en & cacheEntryMemA_line_words_2_MPORT_mask) begin
      cacheEntryMemA_line_words_2[cacheEntryMemA_line_words_2_MPORT_addr] <= cacheEntryMemA_line_words_2_MPORT_data; // @[Cache.scala 115:35]
    end
    cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemA_line_words_3_MPORT_en & cacheEntryMemA_line_words_3_MPORT_mask) begin
      cacheEntryMemA_line_words_3[cacheEntryMemA_line_words_3_MPORT_addr] <= cacheEntryMemA_line_words_3_MPORT_data; // @[Cache.scala 115:35]
    end
    cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemB_valid_MPORT_1_en & cacheEntryMemB_valid_MPORT_1_mask) begin
      cacheEntryMemB_valid[cacheEntryMemB_valid_MPORT_1_addr] <= cacheEntryMemB_valid_MPORT_1_data; // @[Cache.scala 116:35]
    end
    cacheEntryMemB_valid_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_valid_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemB_dirty_MPORT_1_en & cacheEntryMemB_dirty_MPORT_1_mask) begin
      cacheEntryMemB_dirty[cacheEntryMemB_dirty_MPORT_1_addr] <= cacheEntryMemB_dirty_MPORT_1_data; // @[Cache.scala 116:35]
    end
    cacheEntryMemB_dirty_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_dirty_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemB_tag_MPORT_1_en & cacheEntryMemB_tag_MPORT_1_mask) begin
      cacheEntryMemB_tag[cacheEntryMemB_tag_MPORT_1_addr] <= cacheEntryMemB_tag_MPORT_1_data; // @[Cache.scala 116:35]
    end
    cacheEntryMemB_tag_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_tag_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemB_line_words_0_MPORT_1_en & cacheEntryMemB_line_words_0_MPORT_1_mask) begin
      cacheEntryMemB_line_words_0[cacheEntryMemB_line_words_0_MPORT_1_addr] <= cacheEntryMemB_line_words_0_MPORT_1_data; // @[Cache.scala 116:35]
    end
    cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemB_line_words_1_MPORT_1_en & cacheEntryMemB_line_words_1_MPORT_1_mask) begin
      cacheEntryMemB_line_words_1[cacheEntryMemB_line_words_1_MPORT_1_addr] <= cacheEntryMemB_line_words_1_MPORT_1_data; // @[Cache.scala 116:35]
    end
    cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemB_line_words_2_MPORT_1_en & cacheEntryMemB_line_words_2_MPORT_1_mask) begin
      cacheEntryMemB_line_words_2[cacheEntryMemB_line_words_2_MPORT_1_addr] <= cacheEntryMemB_line_words_2_MPORT_1_data; // @[Cache.scala 116:35]
    end
    cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (cacheEntryMemB_line_words_3_MPORT_1_en & cacheEntryMemB_line_words_3_MPORT_1_mask) begin
      cacheEntryMemB_line_words_3[cacheEntryMemB_line_words_3_MPORT_1_addr] <= cacheEntryMemB_line_words_3_MPORT_1_data; // @[Cache.scala 116:35]
    end
    cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[2];
    end
    if (reset) begin // @[Cache.scala 87:25]
      stateReg <= 4'h0; // @[Cache.scala 87:25]
    end else if (4'h0 == stateReg) begin // @[Cache.scala 221:20]
      if (initCounterWrap) begin // @[Cache.scala 224:29]
        stateReg <= 4'h1; // @[Cache.scala 224:40]
      end else begin
        stateReg <= _GEN_67;
      end
    end else if (4'h1 == stateReg) begin // @[Cache.scala 221:20]
      if (start) begin // @[Cache.scala 229:19]
        stateReg <= 4'h2; // @[Cache.scala 229:30]
      end else begin
        stateReg <= _GEN_67;
      end
    end else if (4'h2 == stateReg) begin // @[Cache.scala 221:20]
      stateReg <= _GEN_92;
    end else begin
      stateReg <= _GEN_106;
    end
    if (start) begin // @[Reg.scala 20:18]
      offsetReg <= offsetReg_offset; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_rd <= io_in_rd; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_wr <= io_in_wr; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_addr_tag <= request_addr_tag; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_addr_index <= request_addr_index; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_addr_offset <= request_addr_offset; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_din <= io_in_din; // @[Reg.scala 20:22]
    end
    if (4'h0 == stateReg) begin // @[Cache.scala 221:20]
      doutReg <= _GEN_61;
    end else if (4'h1 == stateReg) begin // @[Cache.scala 221:20]
      doutReg <= _GEN_61;
    end else if (4'h2 == stateReg) begin // @[Cache.scala 221:20]
      if (hit) begin // @[Cache.scala 234:17]
        doutReg <= _GEN_86;
      end else begin
        doutReg <= _GEN_61;
      end
    end else begin
      doutReg <= _GEN_61;
    end
    if (4'h0 == stateReg) begin // @[Cache.scala 221:20]
      validReg <= _GEN_62;
    end else if (4'h1 == stateReg) begin // @[Cache.scala 221:20]
      validReg <= _GEN_62;
    end else if (4'h2 == stateReg) begin // @[Cache.scala 221:20]
      if (hit) begin // @[Cache.scala 234:17]
        validReg <= _GEN_87;
      end else begin
        validReg <= _GEN_62;
      end
    end else begin
      validReg <= _GEN_62;
    end
    if (!(4'h0 == stateReg)) begin // @[Cache.scala 221:20]
      if (!(4'h1 == stateReg)) begin // @[Cache.scala 221:20]
        if (4'h2 == stateReg) begin // @[Cache.scala 221:20]
          if (hit) begin // @[Cache.scala 234:17]
            lruReg <= _lruReg_T_5; // @[Cache.scala 206:12]
          end else begin
            lruReg <= _GEN_91;
          end
        end
      end
    end
    if (4'h0 == stateReg) begin // @[Cache.scala 221:20]
      wayReg <= _nextWay_T_2; // @[Cache.scala 181:11]
    end else if (4'h1 == stateReg) begin // @[Cache.scala 221:20]
      wayReg <= _nextWay_T_2; // @[Cache.scala 181:11]
    end else if (4'h2 == stateReg) begin // @[Cache.scala 221:20]
      if (hit) begin // @[Cache.scala 234:17]
        wayReg <= ~hitA; // @[Cache.scala 207:13]
      end else begin
        wayReg <= _nextWay_T_2; // @[Cache.scala 181:11]
      end
    end else begin
      wayReg <= _nextWay_T_2; // @[Cache.scala 181:11]
    end
    if (!(stateReg == 4'h7)) begin // @[Cache.scala 193:34]
      cacheEntryReg_valid <= _GEN_54;
    end
    cacheEntryReg_dirty <= stateReg == 4'h7 | _GEN_55; // @[Cache.scala 193:34 195:19]
    if (!(stateReg == 4'h7)) begin // @[Cache.scala 193:34]
      if (burstCounterEnable_fill) begin // @[Cache.scala 184:53]
        cacheEntryReg_tag <= requestReg_addr_tag; // @[Cache.scala 187:19]
      end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
        if (nextWay) begin // @[Cache.scala 124:36]
          cacheEntryReg_tag <= cacheEntryMemB_tag_cacheEntryB_data;
        end else begin
          cacheEntryReg_tag <= cacheEntryMemA_tag_cacheEntryA_data;
        end
      end
    end
    if (stateReg == 4'h7) begin // @[Cache.scala 193:34]
      cacheEntryReg_line_words_0 <= cacheEntryReg_entry_line_words_0; // @[Cache.scala 195:19]
    end else if (burstCounterEnable_fill) begin // @[Cache.scala 184:53]
      if (2'h0 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_0 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[Cache.scala 124:36]
        cacheEntryReg_line_words_0 <= cacheEntryMemB_line_words_0_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_0 <= cacheEntryMemA_line_words_0_cacheEntryA_data;
      end
    end
    if (stateReg == 4'h7) begin // @[Cache.scala 193:34]
      cacheEntryReg_line_words_1 <= cacheEntryReg_entry_line_words_1; // @[Cache.scala 195:19]
    end else if (burstCounterEnable_fill) begin // @[Cache.scala 184:53]
      if (2'h1 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_1 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[Cache.scala 124:36]
        cacheEntryReg_line_words_1 <= cacheEntryMemB_line_words_1_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_1 <= cacheEntryMemA_line_words_1_cacheEntryA_data;
      end
    end
    if (stateReg == 4'h7) begin // @[Cache.scala 193:34]
      cacheEntryReg_line_words_2 <= cacheEntryReg_entry_line_words_2; // @[Cache.scala 195:19]
    end else if (burstCounterEnable_fill) begin // @[Cache.scala 184:53]
      if (2'h2 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_2 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[Cache.scala 124:36]
        cacheEntryReg_line_words_2 <= cacheEntryMemB_line_words_2_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_2 <= cacheEntryMemA_line_words_2_cacheEntryA_data;
      end
    end
    if (stateReg == 4'h7) begin // @[Cache.scala 193:34]
      cacheEntryReg_line_words_3 <= cacheEntryReg_entry_line_words_3; // @[Cache.scala 195:19]
    end else if (burstCounterEnable_fill) begin // @[Cache.scala 184:53]
      if (2'h3 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_3 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[Cache.scala 124:36]
        cacheEntryReg_line_words_3 <= cacheEntryMemB_line_words_3_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_3 <= cacheEntryMemA_line_words_3_cacheEntryA_data;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      initCounter <= 1'h0; // @[Counter.scala 61:40]
    end else if (_T) begin // @[Counter.scala 118:16]
      initCounter <= initCounter + 1'h1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      burstCounter <= 2'h0; // @[Counter.scala 61:40]
    end else if (burstCounterEnable) begin // @[Counter.scala 118:16]
      burstCounter <= _wrap_value_T_3; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemA_valid[initvar] = _RAND_0[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemA_dirty[initvar] = _RAND_3[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemA_tag[initvar] = _RAND_6[3:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemA_line_words_0[initvar] = _RAND_9[15:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemA_line_words_1[initvar] = _RAND_12[15:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemA_line_words_2[initvar] = _RAND_15[15:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemA_line_words_3[initvar] = _RAND_18[15:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemB_valid[initvar] = _RAND_21[0:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemB_dirty[initvar] = _RAND_24[0:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemB_tag[initvar] = _RAND_27[3:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemB_line_words_0[initvar] = _RAND_30[15:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemB_line_words_1[initvar] = _RAND_33[15:0];
  _RAND_36 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemB_line_words_2[initvar] = _RAND_36[15:0];
  _RAND_39 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    cacheEntryMemB_line_words_3[initvar] = _RAND_39[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cacheEntryMemA_valid_cacheEntryA_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cacheEntryMemA_valid_cacheEntryA_addr_pipe_0 = _RAND_2[0:0];
  _RAND_4 = {1{`RANDOM}};
  cacheEntryMemA_dirty_cacheEntryA_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cacheEntryMemA_dirty_cacheEntryA_addr_pipe_0 = _RAND_5[0:0];
  _RAND_7 = {1{`RANDOM}};
  cacheEntryMemA_tag_cacheEntryA_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  cacheEntryMemA_tag_cacheEntryA_addr_pipe_0 = _RAND_8[0:0];
  _RAND_10 = {1{`RANDOM}};
  cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0 = _RAND_11[0:0];
  _RAND_13 = {1{`RANDOM}};
  cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0 = _RAND_14[0:0];
  _RAND_16 = {1{`RANDOM}};
  cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0 = _RAND_17[0:0];
  _RAND_19 = {1{`RANDOM}};
  cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0 = _RAND_20[0:0];
  _RAND_22 = {1{`RANDOM}};
  cacheEntryMemB_valid_cacheEntryB_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  cacheEntryMemB_valid_cacheEntryB_addr_pipe_0 = _RAND_23[0:0];
  _RAND_25 = {1{`RANDOM}};
  cacheEntryMemB_dirty_cacheEntryB_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  cacheEntryMemB_dirty_cacheEntryB_addr_pipe_0 = _RAND_26[0:0];
  _RAND_28 = {1{`RANDOM}};
  cacheEntryMemB_tag_cacheEntryB_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  cacheEntryMemB_tag_cacheEntryB_addr_pipe_0 = _RAND_29[0:0];
  _RAND_31 = {1{`RANDOM}};
  cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0 = _RAND_32[0:0];
  _RAND_34 = {1{`RANDOM}};
  cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0 = _RAND_35[0:0];
  _RAND_37 = {1{`RANDOM}};
  cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0 = _RAND_38[0:0];
  _RAND_40 = {1{`RANDOM}};
  cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  stateReg = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  offsetReg = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  requestReg_rd = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  requestReg_wr = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  requestReg_addr_tag = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  requestReg_addr_index = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  requestReg_addr_offset = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  requestReg_din = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  doutReg = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  validReg = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  lruReg = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  wayReg = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  cacheEntryReg_valid = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  cacheEntryReg_dirty = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  cacheEntryReg_tag = _RAND_56[3:0];
  _RAND_57 = {1{`RANDOM}};
  cacheEntryReg_line_words_0 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  cacheEntryReg_line_words_1 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  cacheEntryReg_line_words_2 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  cacheEntryReg_line_words_3 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  initCounter = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  burstCounter = _RAND_62[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReadCache_1(
  input         clock,
  input         reset,
  input         io_enable,
  input         io_in_rd,
  input  [24:0] io_in_addr,
  output [7:0]  io_in_dout,
  output        io_in_wait_n,
  output        io_in_valid,
  output        io_out_rd,
  output [24:0] io_out_addr,
  input  [15:0] io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
`endif // RANDOMIZE_REG_INIT
  reg  cacheEntryMemA_valid [0:3]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [1:0] cacheEntryMemA_valid_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_MPORT_data; // @[ReadCache.scala 112:35]
  wire [1:0] cacheEntryMemA_valid_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_valid_cacheEntryA_en_pipe_0;
  reg [1:0] cacheEntryMemA_valid_cacheEntryA_addr_pipe_0;
  reg [20:0] cacheEntryMemA_tag [0:3]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_tag_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [1:0] cacheEntryMemA_tag_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [20:0] cacheEntryMemA_tag_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [20:0] cacheEntryMemA_tag_MPORT_data; // @[ReadCache.scala 112:35]
  wire [1:0] cacheEntryMemA_tag_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_tag_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_tag_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_tag_cacheEntryA_en_pipe_0;
  reg [1:0] cacheEntryMemA_tag_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_0 [0:3]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_0_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [1:0] cacheEntryMemA_line_words_0_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_0_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_0_MPORT_data; // @[ReadCache.scala 112:35]
  wire [1:0] cacheEntryMemA_line_words_0_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_0_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_0_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0;
  reg [1:0] cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_1 [0:3]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_1_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [1:0] cacheEntryMemA_line_words_1_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_1_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_1_MPORT_data; // @[ReadCache.scala 112:35]
  wire [1:0] cacheEntryMemA_line_words_1_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_1_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_1_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0;
  reg [1:0] cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_2 [0:3]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_2_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [1:0] cacheEntryMemA_line_words_2_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_2_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_2_MPORT_data; // @[ReadCache.scala 112:35]
  wire [1:0] cacheEntryMemA_line_words_2_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_2_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_2_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0;
  reg [1:0] cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_3 [0:3]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_3_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [1:0] cacheEntryMemA_line_words_3_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_3_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_3_MPORT_data; // @[ReadCache.scala 112:35]
  wire [1:0] cacheEntryMemA_line_words_3_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_3_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_3_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0;
  reg [1:0] cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0;
  reg  cacheEntryMemB_valid [0:3]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [1:0] cacheEntryMemB_valid_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [1:0] cacheEntryMemB_valid_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_valid_cacheEntryB_en_pipe_0;
  reg [1:0] cacheEntryMemB_valid_cacheEntryB_addr_pipe_0;
  reg [20:0] cacheEntryMemB_tag [0:3]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_tag_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [1:0] cacheEntryMemB_tag_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [20:0] cacheEntryMemB_tag_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [20:0] cacheEntryMemB_tag_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [1:0] cacheEntryMemB_tag_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_tag_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_tag_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_tag_cacheEntryB_en_pipe_0;
  reg [1:0] cacheEntryMemB_tag_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_0 [0:3]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_0_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [1:0] cacheEntryMemB_line_words_0_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_0_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_0_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [1:0] cacheEntryMemB_line_words_0_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_0_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_0_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0;
  reg [1:0] cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_1 [0:3]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_1_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [1:0] cacheEntryMemB_line_words_1_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_1_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_1_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [1:0] cacheEntryMemB_line_words_1_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_1_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_1_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0;
  reg [1:0] cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_2 [0:3]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_2_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [1:0] cacheEntryMemB_line_words_2_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_2_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_2_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [1:0] cacheEntryMemB_line_words_2_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_2_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_2_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0;
  reg [1:0] cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_3 [0:3]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_3_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [1:0] cacheEntryMemB_line_words_3_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_3_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_3_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [1:0] cacheEntryMemB_line_words_3_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_3_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_3_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0;
  reg [1:0] cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0;
  reg [2:0] stateReg; // @[ReadCache.scala 84:25]
  wire [2:0] offsetReg_offset = io_in_addr[2:0]; // @[ReadCache.scala 92:22]
  reg [2:0] offsetReg; // @[Reg.scala 19:16]
  wire  _start_T_1 = stateReg == 3'h1; // @[ReadCache.scala 142:48]
  wire  start = io_enable & io_in_rd & stateReg == 3'h1; // @[ReadCache.scala 142:36]
  wire [24:0] _request_WIRE_1 = {{1'd0}, io_in_addr[24:1]};
  wire [1:0] request_addr_offset = _request_WIRE_1[1:0]; // @[Address.scala 78:49]
  wire [1:0] request_addr_index = _request_WIRE_1[3:2]; // @[Address.scala 78:49]
  wire [20:0] request_addr_tag = _request_WIRE_1[24:4]; // @[Address.scala 78:49]
  reg  requestReg_rd; // @[Reg.scala 19:16]
  reg [20:0] requestReg_addr_tag; // @[Reg.scala 19:16]
  reg [1:0] requestReg_addr_index; // @[Reg.scala 19:16]
  reg [1:0] requestReg_addr_offset; // @[Reg.scala 19:16]
  reg [7:0] doutReg; // @[ReadCache.scala 101:20]
  reg  validReg; // @[ReadCache.scala 102:25]
  reg [3:0] lruReg; // @[ReadCache.scala 105:19]
  reg  wayReg; // @[ReadCache.scala 109:23]
  wire [3:0] _nextWay_T = lruReg >> request_addr_index; // @[ReadCache.scala 169:31]
  wire  _nextWay_T_2 = start ? _nextWay_T[0] : wayReg; // @[ReadCache.scala 169:17]
  wire  hitA = cacheEntryMemA_valid_cacheEntryA_data & cacheEntryMemA_tag_cacheEntryA_data == requestReg_addr_tag; // @[Entry.scala 59:42]
  wire  hitB = cacheEntryMemB_valid_cacheEntryB_data & cacheEntryMemB_tag_cacheEntryB_data == requestReg_addr_tag; // @[Entry.scala 59:42]
  wire  hit = hitA | hitB; // @[ReadCache.scala 146:18]
  wire  _GEN_88 = hit ? ~hitA : _nextWay_T_2; // @[ReadCache.scala 169:11 185:13 207:17]
  wire  _GEN_98 = 3'h2 == stateReg ? _GEN_88 : _nextWay_T_2; // @[ReadCache.scala 169:11 194:20]
  wire  _GEN_103 = 3'h1 == stateReg ? _nextWay_T_2 : _GEN_98; // @[ReadCache.scala 169:11 194:20]
  wire  nextWay = 3'h0 == stateReg ? _nextWay_T_2 : _GEN_103; // @[ReadCache.scala 169:11 194:20]
  wire  _cacheEntryReg_T_valid = nextWay ? cacheEntryMemB_valid_cacheEntryB_data : cacheEntryMemA_valid_cacheEntryA_data
    ; // @[ReadCache.scala 121:36]
  wire  _cacheEntryReg_T_1 = stateReg == 3'h2; // @[ReadCache.scala 121:82]
  reg  cacheEntryReg_valid; // @[Reg.scala 19:16]
  reg [20:0] cacheEntryReg_tag; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_0; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_1; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_2; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_3; // @[Reg.scala 19:16]
  wire  _GEN_10 = _cacheEntryReg_T_1 ? _cacheEntryReg_T_valid : cacheEntryReg_valid; // @[Reg.scala 19:16 20:{18,22}]
  wire  _nextCacheEntry_T = stateReg == 3'h5; // @[ReadCache.scala 124:37]
  wire  _T = stateReg == 3'h0; // @[ReadCache.scala 126:17]
  wire  _T_2 = ~wayReg; // @[ReadCache.scala 126:64]
  wire  _T_3 = _nextCacheEntry_T & ~wayReg; // @[ReadCache.scala 126:61]
  wire  _T_7 = _nextCacheEntry_T & wayReg; // @[ReadCache.scala 130:61]
  wire  burstCounterEnable = stateReg == 3'h4 & io_out_valid; // @[ReadCache.scala 135:56]
  reg [1:0] initCounter; // @[Counter.scala 61:40]
  wire  wrap_wrap = initCounter == 2'h3; // @[Counter.scala 73:24]
  wire [1:0] _wrap_value_T_1 = initCounter + 2'h1; // @[Counter.scala 77:24]
  wire  initCounterWrap = _T & wrap_wrap; // @[Counter.scala 118:{16,23}]
  reg [1:0] burstCounter; // @[Counter.scala 61:40]
  wire  wrap_wrap_1 = burstCounter == 2'h3; // @[Counter.scala 73:24]
  wire [1:0] _wrap_value_T_3 = burstCounter + 2'h1; // @[Counter.scala 77:24]
  wire  burstCounterWrap = burstCounterEnable & wrap_wrap_1; // @[Counter.scala 118:{16,23}]
  wire  miss = ~hit; // @[ReadCache.scala 147:14]
  wire  wordDone = burstCounter == 2'h0; // @[ReadCache.scala 153:18]
  wire [24:0] _outAddr_T = {requestReg_addr_tag,requestReg_addr_index,requestReg_addr_offset}; // @[ReadCache.scala 165:11]
  wire [25:0] outAddr = {_outAddr_T, 1'h0}; // @[ReadCache.scala 165:18]
  wire [1:0] n = requestReg_addr_offset + burstCounter; // @[ReadCache.scala 173:57]
  wire [15:0] entry_line_words_0 = 2'h0 == n ? io_out_dout : cacheEntryReg_line_words_0; // @[Entry.scala 92:11 93:{30,30}]
  wire [15:0] entry_line_words_1 = 2'h1 == n ? io_out_dout : cacheEntryReg_line_words_1; // @[Entry.scala 92:11 93:{30,30}]
  wire [15:0] entry_line_words_2 = 2'h2 == n ? io_out_dout : cacheEntryReg_line_words_2; // @[Entry.scala 92:11 93:{30,30}]
  wire [15:0] entry_line_words_3 = 2'h3 == n ? io_out_dout : cacheEntryReg_line_words_3; // @[Entry.scala 92:11 93:{30,30}]
  wire [63:0] _doutReg_ws_T = {entry_line_words_3,entry_line_words_2,entry_line_words_1,entry_line_words_0}; // @[Line.scala 77:32]
  wire [7:0] doutReg_ws_0 = _doutReg_ws_T[7:0]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_1 = _doutReg_ws_T[15:8]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_2 = _doutReg_ws_T[23:16]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_3 = _doutReg_ws_T[31:24]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_4 = _doutReg_ws_T[39:32]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_5 = _doutReg_ws_T[47:40]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_6 = _doutReg_ws_T[55:48]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_7 = _doutReg_ws_T[63:56]; // @[Util.scala 104:11]
  wire [7:0] _GEN_48 = 3'h1 == offsetReg ? doutReg_ws_1 : doutReg_ws_0; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_49 = 3'h2 == offsetReg ? doutReg_ws_2 : _GEN_48; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_50 = 3'h3 == offsetReg ? doutReg_ws_3 : _GEN_49; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_51 = 3'h4 == offsetReg ? doutReg_ws_4 : _GEN_50; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_52 = 3'h5 == offsetReg ? doutReg_ws_5 : _GEN_51; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_53 = 3'h6 == offsetReg ? doutReg_ws_6 : _GEN_52; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_54 = 3'h7 == offsetReg ? doutReg_ws_7 : _GEN_53; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_62 = burstCounterEnable ? _GEN_54 : doutReg; // @[ReadCache.scala 172:53 176:13 101:20]
  wire  _GEN_63 = burstCounterEnable & (requestReg_rd & wordDone); // @[ReadCache.scala 172:53 177:14 102:25]
  wire [63:0] _doutReg_ws_T_1 = {cacheEntryMemA_line_words_3_cacheEntryA_data,
    cacheEntryMemA_line_words_2_cacheEntryA_data,cacheEntryMemA_line_words_1_cacheEntryA_data,
    cacheEntryMemA_line_words_0_cacheEntryA_data}; // @[Line.scala 77:32]
  wire [7:0] doutReg_ws_0_1 = _doutReg_ws_T_1[7:0]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_1_1 = _doutReg_ws_T_1[15:8]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_2_1 = _doutReg_ws_T_1[23:16]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_3_1 = _doutReg_ws_T_1[31:24]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_4_1 = _doutReg_ws_T_1[39:32]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_5_1 = _doutReg_ws_T_1[47:40]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_6_1 = _doutReg_ws_T_1[55:48]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_7_1 = _doutReg_ws_T_1[63:56]; // @[Util.scala 104:11]
  wire [7:0] _GEN_67 = 3'h1 == offsetReg ? doutReg_ws_1_1 : doutReg_ws_0_1; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_68 = 3'h2 == offsetReg ? doutReg_ws_2_1 : _GEN_67; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_69 = 3'h3 == offsetReg ? doutReg_ws_3_1 : _GEN_68; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_70 = 3'h4 == offsetReg ? doutReg_ws_4_1 : _GEN_69; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_71 = 3'h5 == offsetReg ? doutReg_ws_5_1 : _GEN_70; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_72 = 3'h6 == offsetReg ? doutReg_ws_6_1 : _GEN_71; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_73 = 3'h7 == offsetReg ? doutReg_ws_7_1 : _GEN_72; // @[Util.scala 104:{11,11}]
  wire [63:0] _doutReg_ws_T_2 = {cacheEntryMemB_line_words_3_cacheEntryB_data,
    cacheEntryMemB_line_words_2_cacheEntryB_data,cacheEntryMemB_line_words_1_cacheEntryB_data,
    cacheEntryMemB_line_words_0_cacheEntryB_data}; // @[Line.scala 77:32]
  wire [7:0] doutReg_ws_0_2 = _doutReg_ws_T_2[7:0]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_1_2 = _doutReg_ws_T_2[15:8]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_2_2 = _doutReg_ws_T_2[23:16]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_3_2 = _doutReg_ws_T_2[31:24]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_4_2 = _doutReg_ws_T_2[39:32]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_5_2 = _doutReg_ws_T_2[47:40]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_6_2 = _doutReg_ws_T_2[55:48]; // @[Util.scala 104:11]
  wire [7:0] doutReg_ws_7_2 = _doutReg_ws_T_2[63:56]; // @[Util.scala 104:11]
  wire [7:0] _GEN_75 = 3'h1 == offsetReg ? doutReg_ws_1_2 : doutReg_ws_0_2; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_76 = 3'h2 == offsetReg ? doutReg_ws_2_2 : _GEN_75; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_77 = 3'h3 == offsetReg ? doutReg_ws_3_2 : _GEN_76; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_78 = 3'h4 == offsetReg ? doutReg_ws_4_2 : _GEN_77; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_79 = 3'h5 == offsetReg ? doutReg_ws_5_2 : _GEN_78; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_80 = 3'h6 == offsetReg ? doutReg_ws_6_2 : _GEN_79; // @[Util.scala 104:{11,11}]
  wire [7:0] _GEN_81 = 3'h7 == offsetReg ? doutReg_ws_7_2 : _GEN_80; // @[Util.scala 104:{11,11}]
  wire [7:0] _doutReg_T_3 = hitA ? _GEN_73 : _GEN_81; // @[ReadCache.scala 182:19]
  wire [3:0] _lruReg_T = 4'h1 << requestReg_addr_index; // @[ReadCache.scala 184:28]
  wire [3:0] _lruReg_T_1 = lruReg | _lruReg_T; // @[ReadCache.scala 184:28]
  wire [3:0] _lruReg_T_2 = ~lruReg; // @[ReadCache.scala 184:28]
  wire [3:0] _lruReg_T_3 = _lruReg_T_2 | _lruReg_T; // @[ReadCache.scala 184:28]
  wire [3:0] _lruReg_T_4 = ~_lruReg_T_3; // @[ReadCache.scala 184:28]
  wire [3:0] _lruReg_T_5 = hitA ? _lruReg_T_1 : _lruReg_T_4; // @[ReadCache.scala 184:28]
  wire [3:0] _lruReg_T_12 = _T_2 ? _lruReg_T_1 : _lruReg_T_4; // @[ReadCache.scala 190:28]
  wire [2:0] _GEN_82 = miss ? 3'h3 : stateReg; // @[ReadCache.scala 189:14 207:44 84:25]
  wire [3:0] _GEN_83 = miss ? _lruReg_T_12 : lruReg; // @[ReadCache.scala 190:12 105:19 207:44]
  wire [2:0] _GEN_84 = hit ? 3'h1 : _GEN_82; // @[ReadCache.scala 181:14 207:17]
  wire  _GEN_86 = hit | _GEN_63; // @[ReadCache.scala 183:14 207:17]
  wire [2:0] _GEN_89 = io_out_wait_n ? 3'h4 : stateReg; // @[ReadCache.scala 212:{27,38} 84:25]
  wire [2:0] _GEN_90 = burstCounterWrap ? 3'h5 : stateReg; // @[ReadCache.scala 217:{30,41} 84:25]
  wire [2:0] _GEN_91 = 3'h5 == stateReg ? 3'h1 : stateReg; // @[ReadCache.scala 194:20 221:32 84:25]
  wire [2:0] _GEN_92 = 3'h4 == stateReg ? _GEN_90 : _GEN_91; // @[ReadCache.scala 194:20]
  wire [2:0] _GEN_93 = 3'h3 == stateReg ? _GEN_89 : _GEN_92; // @[ReadCache.scala 194:20]
  assign cacheEntryMemA_valid_cacheEntryA_en = cacheEntryMemA_valid_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_valid_cacheEntryA_addr = cacheEntryMemA_valid_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_valid_cacheEntryA_data = cacheEntryMemA_valid[cacheEntryMemA_valid_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_valid_MPORT_data = _nextCacheEntry_T & cacheEntryReg_valid;
  assign cacheEntryMemA_valid_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_valid_MPORT_mask = 1'h1;
  assign cacheEntryMemA_valid_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_tag_cacheEntryA_en = cacheEntryMemA_tag_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_tag_cacheEntryA_addr = cacheEntryMemA_tag_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_tag_cacheEntryA_data = cacheEntryMemA_tag[cacheEntryMemA_tag_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_tag_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_tag : 21'h0;
  assign cacheEntryMemA_tag_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_tag_MPORT_mask = 1'h1;
  assign cacheEntryMemA_tag_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_0_cacheEntryA_en = cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_0_cacheEntryA_addr = cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_0_cacheEntryA_data =
    cacheEntryMemA_line_words_0[cacheEntryMemA_line_words_0_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_line_words_0_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_0 : 16'h0;
  assign cacheEntryMemA_line_words_0_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_0_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_0_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_1_cacheEntryA_en = cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_1_cacheEntryA_addr = cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_1_cacheEntryA_data =
    cacheEntryMemA_line_words_1[cacheEntryMemA_line_words_1_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_line_words_1_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_1 : 16'h0;
  assign cacheEntryMemA_line_words_1_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_1_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_1_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_2_cacheEntryA_en = cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_2_cacheEntryA_addr = cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_2_cacheEntryA_data =
    cacheEntryMemA_line_words_2[cacheEntryMemA_line_words_2_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_line_words_2_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_2 : 16'h0;
  assign cacheEntryMemA_line_words_2_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_2_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_2_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_3_cacheEntryA_en = cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_3_cacheEntryA_addr = cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_3_cacheEntryA_data =
    cacheEntryMemA_line_words_3[cacheEntryMemA_line_words_3_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_line_words_3_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_3 : 16'h0;
  assign cacheEntryMemA_line_words_3_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_3_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_3_MPORT_en = _T | _T_3;
  assign cacheEntryMemB_valid_cacheEntryB_en = cacheEntryMemB_valid_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_valid_cacheEntryB_addr = cacheEntryMemB_valid_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_valid_cacheEntryB_data = cacheEntryMemB_valid[cacheEntryMemB_valid_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_valid_MPORT_1_data = _nextCacheEntry_T & cacheEntryReg_valid;
  assign cacheEntryMemB_valid_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_valid_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_valid_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_tag_cacheEntryB_en = cacheEntryMemB_tag_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_tag_cacheEntryB_addr = cacheEntryMemB_tag_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_tag_cacheEntryB_data = cacheEntryMemB_tag[cacheEntryMemB_tag_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_tag_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_tag : 21'h0;
  assign cacheEntryMemB_tag_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_tag_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_tag_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_0_cacheEntryB_en = cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_0_cacheEntryB_addr = cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_0_cacheEntryB_data =
    cacheEntryMemB_line_words_0[cacheEntryMemB_line_words_0_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_line_words_0_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_0 : 16'h0;
  assign cacheEntryMemB_line_words_0_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_0_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_0_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_1_cacheEntryB_en = cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_1_cacheEntryB_addr = cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_1_cacheEntryB_data =
    cacheEntryMemB_line_words_1[cacheEntryMemB_line_words_1_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_line_words_1_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_1 : 16'h0;
  assign cacheEntryMemB_line_words_1_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_1_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_1_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_2_cacheEntryB_en = cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_2_cacheEntryB_addr = cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_2_cacheEntryB_data =
    cacheEntryMemB_line_words_2[cacheEntryMemB_line_words_2_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_line_words_2_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_2 : 16'h0;
  assign cacheEntryMemB_line_words_2_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_2_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_2_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_3_cacheEntryB_en = cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_3_cacheEntryB_addr = cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_3_cacheEntryB_data =
    cacheEntryMemB_line_words_3[cacheEntryMemB_line_words_3_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_line_words_3_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_3 : 16'h0;
  assign cacheEntryMemB_line_words_3_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_3_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_3_MPORT_1_en = _T | _T_7;
  assign io_in_dout = doutReg; // @[ReadCache.scala 227:14]
  assign io_in_wait_n = io_enable & _start_T_1; // @[ReadCache.scala 143:26]
  assign io_in_valid = validReg; // @[ReadCache.scala 226:15]
  assign io_out_rd = stateReg == 3'h3; // @[ReadCache.scala 228:25]
  assign io_out_addr = outAddr[24:0]; // @[ReadCache.scala 230:15]
  always @(posedge clock) begin
    if (cacheEntryMemA_valid_MPORT_en & cacheEntryMemA_valid_MPORT_mask) begin
      cacheEntryMemA_valid[cacheEntryMemA_valid_MPORT_addr] <= cacheEntryMemA_valid_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_valid_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_valid_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[3:2];
    end
    if (cacheEntryMemA_tag_MPORT_en & cacheEntryMemA_tag_MPORT_mask) begin
      cacheEntryMemA_tag[cacheEntryMemA_tag_MPORT_addr] <= cacheEntryMemA_tag_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_tag_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_tag_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[3:2];
    end
    if (cacheEntryMemA_line_words_0_MPORT_en & cacheEntryMemA_line_words_0_MPORT_mask) begin
      cacheEntryMemA_line_words_0[cacheEntryMemA_line_words_0_MPORT_addr] <= cacheEntryMemA_line_words_0_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[3:2];
    end
    if (cacheEntryMemA_line_words_1_MPORT_en & cacheEntryMemA_line_words_1_MPORT_mask) begin
      cacheEntryMemA_line_words_1[cacheEntryMemA_line_words_1_MPORT_addr] <= cacheEntryMemA_line_words_1_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[3:2];
    end
    if (cacheEntryMemA_line_words_2_MPORT_en & cacheEntryMemA_line_words_2_MPORT_mask) begin
      cacheEntryMemA_line_words_2[cacheEntryMemA_line_words_2_MPORT_addr] <= cacheEntryMemA_line_words_2_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[3:2];
    end
    if (cacheEntryMemA_line_words_3_MPORT_en & cacheEntryMemA_line_words_3_MPORT_mask) begin
      cacheEntryMemA_line_words_3[cacheEntryMemA_line_words_3_MPORT_addr] <= cacheEntryMemA_line_words_3_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[3:2];
    end
    if (cacheEntryMemB_valid_MPORT_1_en & cacheEntryMemB_valid_MPORT_1_mask) begin
      cacheEntryMemB_valid[cacheEntryMemB_valid_MPORT_1_addr] <= cacheEntryMemB_valid_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_valid_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_valid_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[3:2];
    end
    if (cacheEntryMemB_tag_MPORT_1_en & cacheEntryMemB_tag_MPORT_1_mask) begin
      cacheEntryMemB_tag[cacheEntryMemB_tag_MPORT_1_addr] <= cacheEntryMemB_tag_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_tag_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_tag_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[3:2];
    end
    if (cacheEntryMemB_line_words_0_MPORT_1_en & cacheEntryMemB_line_words_0_MPORT_1_mask) begin
      cacheEntryMemB_line_words_0[cacheEntryMemB_line_words_0_MPORT_1_addr] <= cacheEntryMemB_line_words_0_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[3:2];
    end
    if (cacheEntryMemB_line_words_1_MPORT_1_en & cacheEntryMemB_line_words_1_MPORT_1_mask) begin
      cacheEntryMemB_line_words_1[cacheEntryMemB_line_words_1_MPORT_1_addr] <= cacheEntryMemB_line_words_1_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[3:2];
    end
    if (cacheEntryMemB_line_words_2_MPORT_1_en & cacheEntryMemB_line_words_2_MPORT_1_mask) begin
      cacheEntryMemB_line_words_2[cacheEntryMemB_line_words_2_MPORT_1_addr] <= cacheEntryMemB_line_words_2_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[3:2];
    end
    if (cacheEntryMemB_line_words_3_MPORT_1_en & cacheEntryMemB_line_words_3_MPORT_1_mask) begin
      cacheEntryMemB_line_words_3[cacheEntryMemB_line_words_3_MPORT_1_addr] <= cacheEntryMemB_line_words_3_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[3:2];
    end
    if (reset) begin // @[ReadCache.scala 84:25]
      stateReg <= 3'h0; // @[ReadCache.scala 84:25]
    end else if (3'h0 == stateReg) begin // @[ReadCache.scala 194:20]
      if (initCounterWrap) begin // @[ReadCache.scala 197:29]
        stateReg <= 3'h1; // @[ReadCache.scala 197:40]
      end
    end else if (3'h1 == stateReg) begin // @[ReadCache.scala 194:20]
      if (start) begin // @[ReadCache.scala 202:19]
        stateReg <= 3'h2; // @[ReadCache.scala 202:30]
      end
    end else if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
      stateReg <= _GEN_84;
    end else begin
      stateReg <= _GEN_93;
    end
    if (start) begin // @[Reg.scala 20:18]
      offsetReg <= offsetReg_offset; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_rd <= io_in_rd; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_addr_tag <= request_addr_tag; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_addr_index <= request_addr_index; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_addr_offset <= request_addr_offset; // @[Reg.scala 20:22]
    end
    if (3'h0 == stateReg) begin // @[ReadCache.scala 194:20]
      doutReg <= _GEN_62;
    end else if (3'h1 == stateReg) begin // @[ReadCache.scala 194:20]
      doutReg <= _GEN_62;
    end else if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
      if (hit) begin // @[ReadCache.scala 207:17]
        doutReg <= _doutReg_T_3; // @[ReadCache.scala 182:13]
      end else begin
        doutReg <= _GEN_62;
      end
    end else begin
      doutReg <= _GEN_62;
    end
    if (3'h0 == stateReg) begin // @[ReadCache.scala 194:20]
      validReg <= _GEN_63;
    end else if (3'h1 == stateReg) begin // @[ReadCache.scala 194:20]
      validReg <= _GEN_63;
    end else if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
      validReg <= _GEN_86;
    end else begin
      validReg <= _GEN_63;
    end
    if (!(3'h0 == stateReg)) begin // @[ReadCache.scala 194:20]
      if (!(3'h1 == stateReg)) begin // @[ReadCache.scala 194:20]
        if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
          if (hit) begin // @[ReadCache.scala 207:17]
            lruReg <= _lruReg_T_5; // @[ReadCache.scala 184:12]
          end else begin
            lruReg <= _GEN_83;
          end
        end
      end
    end
    if (3'h0 == stateReg) begin // @[ReadCache.scala 194:20]
      wayReg <= _nextWay_T_2; // @[ReadCache.scala 169:11]
    end else if (3'h1 == stateReg) begin // @[ReadCache.scala 194:20]
      wayReg <= _nextWay_T_2; // @[ReadCache.scala 169:11]
    end else if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
      if (hit) begin // @[ReadCache.scala 207:17]
        wayReg <= ~hitA; // @[ReadCache.scala 185:13]
      end else begin
        wayReg <= _nextWay_T_2; // @[ReadCache.scala 169:11]
      end
    end else begin
      wayReg <= _nextWay_T_2; // @[ReadCache.scala 169:11]
    end
    cacheEntryReg_valid <= burstCounterEnable | _GEN_10; // @[ReadCache.scala 172:53 175:19]
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      cacheEntryReg_tag <= requestReg_addr_tag; // @[ReadCache.scala 175:19]
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_tag <= cacheEntryMemB_tag_cacheEntryB_data;
      end else begin
        cacheEntryReg_tag <= cacheEntryMemA_tag_cacheEntryA_data;
      end
    end
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      if (2'h0 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_0 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_line_words_0 <= cacheEntryMemB_line_words_0_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_0 <= cacheEntryMemA_line_words_0_cacheEntryA_data;
      end
    end
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      if (2'h1 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_1 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_line_words_1 <= cacheEntryMemB_line_words_1_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_1 <= cacheEntryMemA_line_words_1_cacheEntryA_data;
      end
    end
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      if (2'h2 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_2 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_line_words_2 <= cacheEntryMemB_line_words_2_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_2 <= cacheEntryMemA_line_words_2_cacheEntryA_data;
      end
    end
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      if (2'h3 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_3 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_line_words_3 <= cacheEntryMemB_line_words_3_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_3 <= cacheEntryMemA_line_words_3_cacheEntryA_data;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      initCounter <= 2'h0; // @[Counter.scala 61:40]
    end else if (_T) begin // @[Counter.scala 118:16]
      initCounter <= _wrap_value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      burstCounter <= 2'h0; // @[Counter.scala 61:40]
    end else if (burstCounterEnable) begin // @[Counter.scala 118:16]
      burstCounter <= _wrap_value_T_3; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    cacheEntryMemA_valid[initvar] = _RAND_0[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    cacheEntryMemA_tag[initvar] = _RAND_3[20:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    cacheEntryMemA_line_words_0[initvar] = _RAND_6[15:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    cacheEntryMemA_line_words_1[initvar] = _RAND_9[15:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    cacheEntryMemA_line_words_2[initvar] = _RAND_12[15:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    cacheEntryMemA_line_words_3[initvar] = _RAND_15[15:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    cacheEntryMemB_valid[initvar] = _RAND_18[0:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    cacheEntryMemB_tag[initvar] = _RAND_21[20:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    cacheEntryMemB_line_words_0[initvar] = _RAND_24[15:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    cacheEntryMemB_line_words_1[initvar] = _RAND_27[15:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    cacheEntryMemB_line_words_2[initvar] = _RAND_30[15:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    cacheEntryMemB_line_words_3[initvar] = _RAND_33[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cacheEntryMemA_valid_cacheEntryA_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cacheEntryMemA_valid_cacheEntryA_addr_pipe_0 = _RAND_2[1:0];
  _RAND_4 = {1{`RANDOM}};
  cacheEntryMemA_tag_cacheEntryA_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cacheEntryMemA_tag_cacheEntryA_addr_pipe_0 = _RAND_5[1:0];
  _RAND_7 = {1{`RANDOM}};
  cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0 = _RAND_8[1:0];
  _RAND_10 = {1{`RANDOM}};
  cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0 = _RAND_11[1:0];
  _RAND_13 = {1{`RANDOM}};
  cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0 = _RAND_14[1:0];
  _RAND_16 = {1{`RANDOM}};
  cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0 = _RAND_17[1:0];
  _RAND_19 = {1{`RANDOM}};
  cacheEntryMemB_valid_cacheEntryB_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  cacheEntryMemB_valid_cacheEntryB_addr_pipe_0 = _RAND_20[1:0];
  _RAND_22 = {1{`RANDOM}};
  cacheEntryMemB_tag_cacheEntryB_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  cacheEntryMemB_tag_cacheEntryB_addr_pipe_0 = _RAND_23[1:0];
  _RAND_25 = {1{`RANDOM}};
  cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0 = _RAND_26[1:0];
  _RAND_28 = {1{`RANDOM}};
  cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0 = _RAND_29[1:0];
  _RAND_31 = {1{`RANDOM}};
  cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0 = _RAND_32[1:0];
  _RAND_34 = {1{`RANDOM}};
  cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  stateReg = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  offsetReg = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  requestReg_rd = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  requestReg_addr_tag = _RAND_39[20:0];
  _RAND_40 = {1{`RANDOM}};
  requestReg_addr_index = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  requestReg_addr_offset = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  doutReg = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  validReg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  lruReg = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  wayReg = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  cacheEntryReg_valid = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  cacheEntryReg_tag = _RAND_47[20:0];
  _RAND_48 = {1{`RANDOM}};
  cacheEntryReg_line_words_0 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  cacheEntryReg_line_words_1 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  cacheEntryReg_line_words_2 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  cacheEntryReg_line_words_3 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  initCounter = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  burstCounter = _RAND_53[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReadCache_3(
  input         clock,
  input         reset,
  input         io_enable,
  input         io_in_rd,
  input  [31:0] io_in_addr,
  output [63:0] io_in_dout,
  output        io_in_wait_n,
  output        io_in_valid,
  output        io_out_rd,
  output [24:0] io_out_addr,
  input  [15:0] io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
`endif // RANDOMIZE_REG_INIT
  reg  cacheEntryMemA_valid [0:7]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [2:0] cacheEntryMemA_valid_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_MPORT_data; // @[ReadCache.scala 112:35]
  wire [2:0] cacheEntryMemA_valid_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_valid_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_valid_cacheEntryA_en_pipe_0;
  reg [2:0] cacheEntryMemA_valid_cacheEntryA_addr_pipe_0;
  reg [26:0] cacheEntryMemA_tag [0:7]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_tag_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [2:0] cacheEntryMemA_tag_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [26:0] cacheEntryMemA_tag_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [26:0] cacheEntryMemA_tag_MPORT_data; // @[ReadCache.scala 112:35]
  wire [2:0] cacheEntryMemA_tag_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_tag_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_tag_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_tag_cacheEntryA_en_pipe_0;
  reg [2:0] cacheEntryMemA_tag_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_0 [0:7]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_0_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [2:0] cacheEntryMemA_line_words_0_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_0_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_0_MPORT_data; // @[ReadCache.scala 112:35]
  wire [2:0] cacheEntryMemA_line_words_0_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_0_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_0_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0;
  reg [2:0] cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_1 [0:7]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_1_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [2:0] cacheEntryMemA_line_words_1_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_1_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_1_MPORT_data; // @[ReadCache.scala 112:35]
  wire [2:0] cacheEntryMemA_line_words_1_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_1_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_1_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0;
  reg [2:0] cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_2 [0:7]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_2_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [2:0] cacheEntryMemA_line_words_2_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_2_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_2_MPORT_data; // @[ReadCache.scala 112:35]
  wire [2:0] cacheEntryMemA_line_words_2_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_2_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_2_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0;
  reg [2:0] cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0;
  reg [15:0] cacheEntryMemA_line_words_3 [0:7]; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_3_cacheEntryA_en; // @[ReadCache.scala 112:35]
  wire [2:0] cacheEntryMemA_line_words_3_cacheEntryA_addr; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_3_cacheEntryA_data; // @[ReadCache.scala 112:35]
  wire [15:0] cacheEntryMemA_line_words_3_MPORT_data; // @[ReadCache.scala 112:35]
  wire [2:0] cacheEntryMemA_line_words_3_MPORT_addr; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_3_MPORT_mask; // @[ReadCache.scala 112:35]
  wire  cacheEntryMemA_line_words_3_MPORT_en; // @[ReadCache.scala 112:35]
  reg  cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0;
  reg [2:0] cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0;
  reg  cacheEntryMemB_valid [0:7]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [2:0] cacheEntryMemB_valid_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [2:0] cacheEntryMemB_valid_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_valid_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_valid_cacheEntryB_en_pipe_0;
  reg [2:0] cacheEntryMemB_valid_cacheEntryB_addr_pipe_0;
  reg [26:0] cacheEntryMemB_tag [0:7]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_tag_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [2:0] cacheEntryMemB_tag_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [26:0] cacheEntryMemB_tag_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [26:0] cacheEntryMemB_tag_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [2:0] cacheEntryMemB_tag_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_tag_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_tag_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_tag_cacheEntryB_en_pipe_0;
  reg [2:0] cacheEntryMemB_tag_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_0 [0:7]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_0_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [2:0] cacheEntryMemB_line_words_0_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_0_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_0_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [2:0] cacheEntryMemB_line_words_0_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_0_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_0_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0;
  reg [2:0] cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_1 [0:7]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_1_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [2:0] cacheEntryMemB_line_words_1_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_1_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_1_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [2:0] cacheEntryMemB_line_words_1_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_1_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_1_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0;
  reg [2:0] cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_2 [0:7]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_2_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [2:0] cacheEntryMemB_line_words_2_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_2_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_2_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [2:0] cacheEntryMemB_line_words_2_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_2_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_2_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0;
  reg [2:0] cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0;
  reg [15:0] cacheEntryMemB_line_words_3 [0:7]; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_3_cacheEntryB_en; // @[ReadCache.scala 113:35]
  wire [2:0] cacheEntryMemB_line_words_3_cacheEntryB_addr; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_3_cacheEntryB_data; // @[ReadCache.scala 113:35]
  wire [15:0] cacheEntryMemB_line_words_3_MPORT_1_data; // @[ReadCache.scala 113:35]
  wire [2:0] cacheEntryMemB_line_words_3_MPORT_1_addr; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_3_MPORT_1_mask; // @[ReadCache.scala 113:35]
  wire  cacheEntryMemB_line_words_3_MPORT_1_en; // @[ReadCache.scala 113:35]
  reg  cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0;
  reg [2:0] cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0;
  reg [2:0] stateReg; // @[ReadCache.scala 84:25]
  wire  _start_T_1 = stateReg == 3'h1; // @[ReadCache.scala 142:48]
  wire  start = io_enable & io_in_rd & stateReg == 3'h1; // @[ReadCache.scala 142:36]
  wire [31:0] _request_WIRE_1 = {{1'd0}, io_in_addr[31:1]};
  wire [1:0] request_addr_offset = _request_WIRE_1[1:0]; // @[Address.scala 78:49]
  wire [2:0] request_addr_index = _request_WIRE_1[4:2]; // @[Address.scala 78:49]
  wire [26:0] request_addr_tag = _request_WIRE_1[31:5]; // @[Address.scala 78:49]
  reg  requestReg_rd; // @[Reg.scala 19:16]
  reg [26:0] requestReg_addr_tag; // @[Reg.scala 19:16]
  reg [2:0] requestReg_addr_index; // @[Reg.scala 19:16]
  reg [1:0] requestReg_addr_offset; // @[Reg.scala 19:16]
  reg [63:0] doutReg; // @[ReadCache.scala 101:20]
  reg  validReg; // @[ReadCache.scala 102:25]
  reg [7:0] lruReg; // @[ReadCache.scala 105:19]
  reg  wayReg; // @[ReadCache.scala 109:23]
  wire [7:0] _nextWay_T = lruReg >> request_addr_index; // @[ReadCache.scala 169:31]
  wire  _nextWay_T_2 = start ? _nextWay_T[0] : wayReg; // @[ReadCache.scala 169:17]
  wire  hitA = cacheEntryMemA_valid_cacheEntryA_data & cacheEntryMemA_tag_cacheEntryA_data == requestReg_addr_tag; // @[Entry.scala 59:42]
  wire  hitB = cacheEntryMemB_valid_cacheEntryB_data & cacheEntryMemB_tag_cacheEntryB_data == requestReg_addr_tag; // @[Entry.scala 59:42]
  wire  hit = hitA | hitB; // @[ReadCache.scala 146:18]
  wire  _GEN_64 = hit ? ~hitA : _nextWay_T_2; // @[ReadCache.scala 169:11 185:13 207:17]
  wire  _GEN_74 = 3'h2 == stateReg ? _GEN_64 : _nextWay_T_2; // @[ReadCache.scala 169:11 194:20]
  wire  _GEN_79 = 3'h1 == stateReg ? _nextWay_T_2 : _GEN_74; // @[ReadCache.scala 169:11 194:20]
  wire  nextWay = 3'h0 == stateReg ? _nextWay_T_2 : _GEN_79; // @[ReadCache.scala 169:11 194:20]
  wire  _cacheEntryReg_T_valid = nextWay ? cacheEntryMemB_valid_cacheEntryB_data : cacheEntryMemA_valid_cacheEntryA_data
    ; // @[ReadCache.scala 121:36]
  wire  _cacheEntryReg_T_1 = stateReg == 3'h2; // @[ReadCache.scala 121:82]
  reg  cacheEntryReg_valid; // @[Reg.scala 19:16]
  reg [26:0] cacheEntryReg_tag; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_0; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_1; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_2; // @[Reg.scala 19:16]
  reg [15:0] cacheEntryReg_line_words_3; // @[Reg.scala 19:16]
  wire  _GEN_10 = _cacheEntryReg_T_1 ? _cacheEntryReg_T_valid : cacheEntryReg_valid; // @[Reg.scala 19:16 20:{18,22}]
  wire  _nextCacheEntry_T = stateReg == 3'h5; // @[ReadCache.scala 124:37]
  wire  _T = stateReg == 3'h0; // @[ReadCache.scala 126:17]
  wire  _T_2 = ~wayReg; // @[ReadCache.scala 126:64]
  wire  _T_3 = _nextCacheEntry_T & ~wayReg; // @[ReadCache.scala 126:61]
  wire  _T_7 = _nextCacheEntry_T & wayReg; // @[ReadCache.scala 130:61]
  wire  burstCounterEnable = stateReg == 3'h4 & io_out_valid; // @[ReadCache.scala 135:56]
  reg [2:0] initCounter; // @[Counter.scala 61:40]
  wire  wrap_wrap = initCounter == 3'h7; // @[Counter.scala 73:24]
  wire [2:0] _wrap_value_T_1 = initCounter + 3'h1; // @[Counter.scala 77:24]
  wire  initCounterWrap = _T & wrap_wrap; // @[Counter.scala 118:{16,23}]
  reg [1:0] burstCounter; // @[Counter.scala 61:40]
  wire  wrap_wrap_1 = burstCounter == 2'h3; // @[Counter.scala 73:24]
  wire [1:0] _wrap_value_T_3 = burstCounter + 2'h1; // @[Counter.scala 77:24]
  wire  burstCounterWrap = burstCounterEnable & wrap_wrap_1; // @[Counter.scala 118:{16,23}]
  wire  miss = ~hit; // @[ReadCache.scala 147:14]
  wire [31:0] _outAddr_T = {requestReg_addr_tag,requestReg_addr_index,requestReg_addr_offset}; // @[ReadCache.scala 165:11]
  wire [32:0] outAddr = {_outAddr_T, 1'h0}; // @[ReadCache.scala 165:18]
  wire [1:0] n = requestReg_addr_offset + burstCounter; // @[ReadCache.scala 173:57]
  wire [15:0] entry_line_words_0 = 2'h0 == n ? io_out_dout : cacheEntryReg_line_words_0; // @[Entry.scala 92:11 93:{30,30}]
  wire [15:0] entry_line_words_1 = 2'h1 == n ? io_out_dout : cacheEntryReg_line_words_1; // @[Entry.scala 92:11 93:{30,30}]
  wire [15:0] entry_line_words_2 = 2'h2 == n ? io_out_dout : cacheEntryReg_line_words_2; // @[Entry.scala 92:11 93:{30,30}]
  wire [15:0] entry_line_words_3 = 2'h3 == n ? io_out_dout : cacheEntryReg_line_words_3; // @[Entry.scala 92:11 93:{30,30}]
  wire [63:0] doutReg_ws_0 = {entry_line_words_3,entry_line_words_2,entry_line_words_1,entry_line_words_0}; // @[Line.scala 77:32]
  wire [63:0] _doutReg_T_14 = {doutReg_ws_0[7:0],doutReg_ws_0[15:8],doutReg_ws_0[23:16],doutReg_ws_0[31:24],doutReg_ws_0
    [39:32],doutReg_ws_0[47:40],doutReg_ws_0[55:48],doutReg_ws_0[63:56]}; // @[Util.scala 114:49]
  wire [63:0] _GEN_54 = burstCounterEnable ? _doutReg_T_14 : doutReg; // @[ReadCache.scala 172:53 176:13 101:20]
  wire  _GEN_55 = burstCounterEnable & (requestReg_rd & wrap_wrap_1); // @[ReadCache.scala 172:53 177:14 102:25]
  wire [63:0] doutReg_ws_0_1 = {cacheEntryMemA_line_words_3_cacheEntryA_data,
    cacheEntryMemA_line_words_2_cacheEntryA_data,cacheEntryMemA_line_words_1_cacheEntryA_data,
    cacheEntryMemA_line_words_0_cacheEntryA_data}; // @[Line.scala 77:32]
  wire [63:0] _doutReg_T_29 = {doutReg_ws_0_1[7:0],doutReg_ws_0_1[15:8],doutReg_ws_0_1[23:16],doutReg_ws_0_1[31:24],
    doutReg_ws_0_1[39:32],doutReg_ws_0_1[47:40],doutReg_ws_0_1[55:48],doutReg_ws_0_1[63:56]}; // @[Util.scala 114:49]
  wire [63:0] doutReg_ws_0_2 = {cacheEntryMemB_line_words_3_cacheEntryB_data,
    cacheEntryMemB_line_words_2_cacheEntryB_data,cacheEntryMemB_line_words_1_cacheEntryB_data,
    cacheEntryMemB_line_words_0_cacheEntryB_data}; // @[Line.scala 77:32]
  wire [63:0] _doutReg_T_44 = {doutReg_ws_0_2[7:0],doutReg_ws_0_2[15:8],doutReg_ws_0_2[23:16],doutReg_ws_0_2[31:24],
    doutReg_ws_0_2[39:32],doutReg_ws_0_2[47:40],doutReg_ws_0_2[55:48],doutReg_ws_0_2[63:56]}; // @[Util.scala 114:49]
  wire [63:0] _doutReg_T_45 = hitA ? _doutReg_T_29 : _doutReg_T_44; // @[ReadCache.scala 182:19]
  wire [7:0] _lruReg_T = 8'h1 << requestReg_addr_index; // @[ReadCache.scala 184:28]
  wire [7:0] _lruReg_T_1 = lruReg | _lruReg_T; // @[ReadCache.scala 184:28]
  wire [7:0] _lruReg_T_2 = ~lruReg; // @[ReadCache.scala 184:28]
  wire [7:0] _lruReg_T_3 = _lruReg_T_2 | _lruReg_T; // @[ReadCache.scala 184:28]
  wire [7:0] _lruReg_T_4 = ~_lruReg_T_3; // @[ReadCache.scala 184:28]
  wire [7:0] _lruReg_T_5 = hitA ? _lruReg_T_1 : _lruReg_T_4; // @[ReadCache.scala 184:28]
  wire [7:0] _lruReg_T_12 = _T_2 ? _lruReg_T_1 : _lruReg_T_4; // @[ReadCache.scala 190:28]
  wire [2:0] _GEN_58 = miss ? 3'h3 : stateReg; // @[ReadCache.scala 189:14 207:44 84:25]
  wire [7:0] _GEN_59 = miss ? _lruReg_T_12 : lruReg; // @[ReadCache.scala 190:12 105:19 207:44]
  wire [2:0] _GEN_60 = hit ? 3'h1 : _GEN_58; // @[ReadCache.scala 181:14 207:17]
  wire  _GEN_62 = hit | _GEN_55; // @[ReadCache.scala 183:14 207:17]
  wire [2:0] _GEN_65 = io_out_wait_n ? 3'h4 : stateReg; // @[ReadCache.scala 212:{27,38} 84:25]
  wire [2:0] _GEN_66 = burstCounterWrap ? 3'h5 : stateReg; // @[ReadCache.scala 217:{30,41} 84:25]
  wire [2:0] _GEN_67 = 3'h5 == stateReg ? 3'h1 : stateReg; // @[ReadCache.scala 194:20 221:32 84:25]
  wire [2:0] _GEN_68 = 3'h4 == stateReg ? _GEN_66 : _GEN_67; // @[ReadCache.scala 194:20]
  wire [2:0] _GEN_69 = 3'h3 == stateReg ? _GEN_65 : _GEN_68; // @[ReadCache.scala 194:20]
  assign cacheEntryMemA_valid_cacheEntryA_en = cacheEntryMemA_valid_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_valid_cacheEntryA_addr = cacheEntryMemA_valid_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_valid_cacheEntryA_data = cacheEntryMemA_valid[cacheEntryMemA_valid_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_valid_MPORT_data = _nextCacheEntry_T & cacheEntryReg_valid;
  assign cacheEntryMemA_valid_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_valid_MPORT_mask = 1'h1;
  assign cacheEntryMemA_valid_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_tag_cacheEntryA_en = cacheEntryMemA_tag_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_tag_cacheEntryA_addr = cacheEntryMemA_tag_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_tag_cacheEntryA_data = cacheEntryMemA_tag[cacheEntryMemA_tag_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_tag_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_tag : 27'h0;
  assign cacheEntryMemA_tag_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_tag_MPORT_mask = 1'h1;
  assign cacheEntryMemA_tag_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_0_cacheEntryA_en = cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_0_cacheEntryA_addr = cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_0_cacheEntryA_data =
    cacheEntryMemA_line_words_0[cacheEntryMemA_line_words_0_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_line_words_0_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_0 : 16'h0;
  assign cacheEntryMemA_line_words_0_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_0_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_0_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_1_cacheEntryA_en = cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_1_cacheEntryA_addr = cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_1_cacheEntryA_data =
    cacheEntryMemA_line_words_1[cacheEntryMemA_line_words_1_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_line_words_1_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_1 : 16'h0;
  assign cacheEntryMemA_line_words_1_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_1_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_1_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_2_cacheEntryA_en = cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_2_cacheEntryA_addr = cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_2_cacheEntryA_data =
    cacheEntryMemA_line_words_2[cacheEntryMemA_line_words_2_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_line_words_2_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_2 : 16'h0;
  assign cacheEntryMemA_line_words_2_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_2_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_2_MPORT_en = _T | _T_3;
  assign cacheEntryMemA_line_words_3_cacheEntryA_en = cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0;
  assign cacheEntryMemA_line_words_3_cacheEntryA_addr = cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0;
  assign cacheEntryMemA_line_words_3_cacheEntryA_data =
    cacheEntryMemA_line_words_3[cacheEntryMemA_line_words_3_cacheEntryA_addr]; // @[ReadCache.scala 112:35]
  assign cacheEntryMemA_line_words_3_MPORT_data = _nextCacheEntry_T ? cacheEntryReg_line_words_3 : 16'h0;
  assign cacheEntryMemA_line_words_3_MPORT_addr = requestReg_addr_index;
  assign cacheEntryMemA_line_words_3_MPORT_mask = 1'h1;
  assign cacheEntryMemA_line_words_3_MPORT_en = _T | _T_3;
  assign cacheEntryMemB_valid_cacheEntryB_en = cacheEntryMemB_valid_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_valid_cacheEntryB_addr = cacheEntryMemB_valid_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_valid_cacheEntryB_data = cacheEntryMemB_valid[cacheEntryMemB_valid_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_valid_MPORT_1_data = _nextCacheEntry_T & cacheEntryReg_valid;
  assign cacheEntryMemB_valid_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_valid_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_valid_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_tag_cacheEntryB_en = cacheEntryMemB_tag_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_tag_cacheEntryB_addr = cacheEntryMemB_tag_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_tag_cacheEntryB_data = cacheEntryMemB_tag[cacheEntryMemB_tag_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_tag_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_tag : 27'h0;
  assign cacheEntryMemB_tag_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_tag_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_tag_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_0_cacheEntryB_en = cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_0_cacheEntryB_addr = cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_0_cacheEntryB_data =
    cacheEntryMemB_line_words_0[cacheEntryMemB_line_words_0_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_line_words_0_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_0 : 16'h0;
  assign cacheEntryMemB_line_words_0_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_0_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_0_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_1_cacheEntryB_en = cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_1_cacheEntryB_addr = cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_1_cacheEntryB_data =
    cacheEntryMemB_line_words_1[cacheEntryMemB_line_words_1_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_line_words_1_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_1 : 16'h0;
  assign cacheEntryMemB_line_words_1_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_1_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_1_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_2_cacheEntryB_en = cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_2_cacheEntryB_addr = cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_2_cacheEntryB_data =
    cacheEntryMemB_line_words_2[cacheEntryMemB_line_words_2_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_line_words_2_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_2 : 16'h0;
  assign cacheEntryMemB_line_words_2_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_2_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_2_MPORT_1_en = _T | _T_7;
  assign cacheEntryMemB_line_words_3_cacheEntryB_en = cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0;
  assign cacheEntryMemB_line_words_3_cacheEntryB_addr = cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0;
  assign cacheEntryMemB_line_words_3_cacheEntryB_data =
    cacheEntryMemB_line_words_3[cacheEntryMemB_line_words_3_cacheEntryB_addr]; // @[ReadCache.scala 113:35]
  assign cacheEntryMemB_line_words_3_MPORT_1_data = _nextCacheEntry_T ? cacheEntryReg_line_words_3 : 16'h0;
  assign cacheEntryMemB_line_words_3_MPORT_1_addr = requestReg_addr_index;
  assign cacheEntryMemB_line_words_3_MPORT_1_mask = 1'h1;
  assign cacheEntryMemB_line_words_3_MPORT_1_en = _T | _T_7;
  assign io_in_dout = doutReg; // @[ReadCache.scala 227:14]
  assign io_in_wait_n = io_enable & _start_T_1; // @[ReadCache.scala 143:26]
  assign io_in_valid = validReg; // @[ReadCache.scala 226:15]
  assign io_out_rd = stateReg == 3'h3; // @[ReadCache.scala 228:25]
  assign io_out_addr = outAddr[24:0]; // @[ReadCache.scala 230:15]
  always @(posedge clock) begin
    if (cacheEntryMemA_valid_MPORT_en & cacheEntryMemA_valid_MPORT_mask) begin
      cacheEntryMemA_valid[cacheEntryMemA_valid_MPORT_addr] <= cacheEntryMemA_valid_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_valid_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_valid_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[4:2];
    end
    if (cacheEntryMemA_tag_MPORT_en & cacheEntryMemA_tag_MPORT_mask) begin
      cacheEntryMemA_tag[cacheEntryMemA_tag_MPORT_addr] <= cacheEntryMemA_tag_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_tag_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_tag_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[4:2];
    end
    if (cacheEntryMemA_line_words_0_MPORT_en & cacheEntryMemA_line_words_0_MPORT_mask) begin
      cacheEntryMemA_line_words_0[cacheEntryMemA_line_words_0_MPORT_addr] <= cacheEntryMemA_line_words_0_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[4:2];
    end
    if (cacheEntryMemA_line_words_1_MPORT_en & cacheEntryMemA_line_words_1_MPORT_mask) begin
      cacheEntryMemA_line_words_1[cacheEntryMemA_line_words_1_MPORT_addr] <= cacheEntryMemA_line_words_1_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[4:2];
    end
    if (cacheEntryMemA_line_words_2_MPORT_en & cacheEntryMemA_line_words_2_MPORT_mask) begin
      cacheEntryMemA_line_words_2[cacheEntryMemA_line_words_2_MPORT_addr] <= cacheEntryMemA_line_words_2_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[4:2];
    end
    if (cacheEntryMemA_line_words_3_MPORT_en & cacheEntryMemA_line_words_3_MPORT_mask) begin
      cacheEntryMemA_line_words_3[cacheEntryMemA_line_words_3_MPORT_addr] <= cacheEntryMemA_line_words_3_MPORT_data; // @[ReadCache.scala 112:35]
    end
    cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0 <= _request_WIRE_1[4:2];
    end
    if (cacheEntryMemB_valid_MPORT_1_en & cacheEntryMemB_valid_MPORT_1_mask) begin
      cacheEntryMemB_valid[cacheEntryMemB_valid_MPORT_1_addr] <= cacheEntryMemB_valid_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_valid_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_valid_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[4:2];
    end
    if (cacheEntryMemB_tag_MPORT_1_en & cacheEntryMemB_tag_MPORT_1_mask) begin
      cacheEntryMemB_tag[cacheEntryMemB_tag_MPORT_1_addr] <= cacheEntryMemB_tag_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_tag_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_tag_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[4:2];
    end
    if (cacheEntryMemB_line_words_0_MPORT_1_en & cacheEntryMemB_line_words_0_MPORT_1_mask) begin
      cacheEntryMemB_line_words_0[cacheEntryMemB_line_words_0_MPORT_1_addr] <= cacheEntryMemB_line_words_0_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[4:2];
    end
    if (cacheEntryMemB_line_words_1_MPORT_1_en & cacheEntryMemB_line_words_1_MPORT_1_mask) begin
      cacheEntryMemB_line_words_1[cacheEntryMemB_line_words_1_MPORT_1_addr] <= cacheEntryMemB_line_words_1_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[4:2];
    end
    if (cacheEntryMemB_line_words_2_MPORT_1_en & cacheEntryMemB_line_words_2_MPORT_1_mask) begin
      cacheEntryMemB_line_words_2[cacheEntryMemB_line_words_2_MPORT_1_addr] <= cacheEntryMemB_line_words_2_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[4:2];
    end
    if (cacheEntryMemB_line_words_3_MPORT_1_en & cacheEntryMemB_line_words_3_MPORT_1_mask) begin
      cacheEntryMemB_line_words_3[cacheEntryMemB_line_words_3_MPORT_1_addr] <= cacheEntryMemB_line_words_3_MPORT_1_data; // @[ReadCache.scala 113:35]
    end
    cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0 <= _request_WIRE_1[4:2];
    end
    if (reset) begin // @[ReadCache.scala 84:25]
      stateReg <= 3'h0; // @[ReadCache.scala 84:25]
    end else if (3'h0 == stateReg) begin // @[ReadCache.scala 194:20]
      if (initCounterWrap) begin // @[ReadCache.scala 197:29]
        stateReg <= 3'h1; // @[ReadCache.scala 197:40]
      end
    end else if (3'h1 == stateReg) begin // @[ReadCache.scala 194:20]
      if (start) begin // @[ReadCache.scala 202:19]
        stateReg <= 3'h2; // @[ReadCache.scala 202:30]
      end
    end else if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
      stateReg <= _GEN_60;
    end else begin
      stateReg <= _GEN_69;
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_rd <= io_in_rd; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_addr_tag <= request_addr_tag; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_addr_index <= request_addr_index; // @[Reg.scala 20:22]
    end
    if (start) begin // @[Reg.scala 20:18]
      requestReg_addr_offset <= request_addr_offset; // @[Reg.scala 20:22]
    end
    if (3'h0 == stateReg) begin // @[ReadCache.scala 194:20]
      doutReg <= _GEN_54;
    end else if (3'h1 == stateReg) begin // @[ReadCache.scala 194:20]
      doutReg <= _GEN_54;
    end else if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
      if (hit) begin // @[ReadCache.scala 207:17]
        doutReg <= _doutReg_T_45; // @[ReadCache.scala 182:13]
      end else begin
        doutReg <= _GEN_54;
      end
    end else begin
      doutReg <= _GEN_54;
    end
    if (3'h0 == stateReg) begin // @[ReadCache.scala 194:20]
      validReg <= _GEN_55;
    end else if (3'h1 == stateReg) begin // @[ReadCache.scala 194:20]
      validReg <= _GEN_55;
    end else if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
      validReg <= _GEN_62;
    end else begin
      validReg <= _GEN_55;
    end
    if (!(3'h0 == stateReg)) begin // @[ReadCache.scala 194:20]
      if (!(3'h1 == stateReg)) begin // @[ReadCache.scala 194:20]
        if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
          if (hit) begin // @[ReadCache.scala 207:17]
            lruReg <= _lruReg_T_5; // @[ReadCache.scala 184:12]
          end else begin
            lruReg <= _GEN_59;
          end
        end
      end
    end
    if (3'h0 == stateReg) begin // @[ReadCache.scala 194:20]
      wayReg <= _nextWay_T_2; // @[ReadCache.scala 169:11]
    end else if (3'h1 == stateReg) begin // @[ReadCache.scala 194:20]
      wayReg <= _nextWay_T_2; // @[ReadCache.scala 169:11]
    end else if (3'h2 == stateReg) begin // @[ReadCache.scala 194:20]
      if (hit) begin // @[ReadCache.scala 207:17]
        wayReg <= ~hitA; // @[ReadCache.scala 185:13]
      end else begin
        wayReg <= _nextWay_T_2; // @[ReadCache.scala 169:11]
      end
    end else begin
      wayReg <= _nextWay_T_2; // @[ReadCache.scala 169:11]
    end
    cacheEntryReg_valid <= burstCounterEnable | _GEN_10; // @[ReadCache.scala 172:53 175:19]
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      cacheEntryReg_tag <= requestReg_addr_tag; // @[ReadCache.scala 175:19]
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_tag <= cacheEntryMemB_tag_cacheEntryB_data;
      end else begin
        cacheEntryReg_tag <= cacheEntryMemA_tag_cacheEntryA_data;
      end
    end
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      if (2'h0 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_0 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_line_words_0 <= cacheEntryMemB_line_words_0_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_0 <= cacheEntryMemA_line_words_0_cacheEntryA_data;
      end
    end
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      if (2'h1 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_1 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_line_words_1 <= cacheEntryMemB_line_words_1_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_1 <= cacheEntryMemA_line_words_1_cacheEntryA_data;
      end
    end
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      if (2'h2 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_2 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_line_words_2 <= cacheEntryMemB_line_words_2_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_2 <= cacheEntryMemA_line_words_2_cacheEntryA_data;
      end
    end
    if (burstCounterEnable) begin // @[ReadCache.scala 172:53]
      if (2'h3 == n) begin // @[Entry.scala 93:30]
        cacheEntryReg_line_words_3 <= io_out_dout; // @[Entry.scala 93:30]
      end
    end else if (_cacheEntryReg_T_1) begin // @[Reg.scala 20:18]
      if (nextWay) begin // @[ReadCache.scala 121:36]
        cacheEntryReg_line_words_3 <= cacheEntryMemB_line_words_3_cacheEntryB_data;
      end else begin
        cacheEntryReg_line_words_3 <= cacheEntryMemA_line_words_3_cacheEntryA_data;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      initCounter <= 3'h0; // @[Counter.scala 61:40]
    end else if (_T) begin // @[Counter.scala 118:16]
      initCounter <= _wrap_value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      burstCounter <= 2'h0; // @[Counter.scala 61:40]
    end else if (burstCounterEnable) begin // @[Counter.scala 118:16]
      burstCounter <= _wrap_value_T_3; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cacheEntryMemA_valid[initvar] = _RAND_0[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cacheEntryMemA_tag[initvar] = _RAND_3[26:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cacheEntryMemA_line_words_0[initvar] = _RAND_6[15:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cacheEntryMemA_line_words_1[initvar] = _RAND_9[15:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cacheEntryMemA_line_words_2[initvar] = _RAND_12[15:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cacheEntryMemA_line_words_3[initvar] = _RAND_15[15:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cacheEntryMemB_valid[initvar] = _RAND_18[0:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cacheEntryMemB_tag[initvar] = _RAND_21[26:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cacheEntryMemB_line_words_0[initvar] = _RAND_24[15:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cacheEntryMemB_line_words_1[initvar] = _RAND_27[15:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cacheEntryMemB_line_words_2[initvar] = _RAND_30[15:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cacheEntryMemB_line_words_3[initvar] = _RAND_33[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cacheEntryMemA_valid_cacheEntryA_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cacheEntryMemA_valid_cacheEntryA_addr_pipe_0 = _RAND_2[2:0];
  _RAND_4 = {1{`RANDOM}};
  cacheEntryMemA_tag_cacheEntryA_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cacheEntryMemA_tag_cacheEntryA_addr_pipe_0 = _RAND_5[2:0];
  _RAND_7 = {1{`RANDOM}};
  cacheEntryMemA_line_words_0_cacheEntryA_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  cacheEntryMemA_line_words_0_cacheEntryA_addr_pipe_0 = _RAND_8[2:0];
  _RAND_10 = {1{`RANDOM}};
  cacheEntryMemA_line_words_1_cacheEntryA_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cacheEntryMemA_line_words_1_cacheEntryA_addr_pipe_0 = _RAND_11[2:0];
  _RAND_13 = {1{`RANDOM}};
  cacheEntryMemA_line_words_2_cacheEntryA_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  cacheEntryMemA_line_words_2_cacheEntryA_addr_pipe_0 = _RAND_14[2:0];
  _RAND_16 = {1{`RANDOM}};
  cacheEntryMemA_line_words_3_cacheEntryA_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  cacheEntryMemA_line_words_3_cacheEntryA_addr_pipe_0 = _RAND_17[2:0];
  _RAND_19 = {1{`RANDOM}};
  cacheEntryMemB_valid_cacheEntryB_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  cacheEntryMemB_valid_cacheEntryB_addr_pipe_0 = _RAND_20[2:0];
  _RAND_22 = {1{`RANDOM}};
  cacheEntryMemB_tag_cacheEntryB_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  cacheEntryMemB_tag_cacheEntryB_addr_pipe_0 = _RAND_23[2:0];
  _RAND_25 = {1{`RANDOM}};
  cacheEntryMemB_line_words_0_cacheEntryB_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  cacheEntryMemB_line_words_0_cacheEntryB_addr_pipe_0 = _RAND_26[2:0];
  _RAND_28 = {1{`RANDOM}};
  cacheEntryMemB_line_words_1_cacheEntryB_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  cacheEntryMemB_line_words_1_cacheEntryB_addr_pipe_0 = _RAND_29[2:0];
  _RAND_31 = {1{`RANDOM}};
  cacheEntryMemB_line_words_2_cacheEntryB_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  cacheEntryMemB_line_words_2_cacheEntryB_addr_pipe_0 = _RAND_32[2:0];
  _RAND_34 = {1{`RANDOM}};
  cacheEntryMemB_line_words_3_cacheEntryB_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  cacheEntryMemB_line_words_3_cacheEntryB_addr_pipe_0 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  stateReg = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  requestReg_rd = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  requestReg_addr_tag = _RAND_38[26:0];
  _RAND_39 = {1{`RANDOM}};
  requestReg_addr_index = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  requestReg_addr_offset = _RAND_40[1:0];
  _RAND_41 = {2{`RANDOM}};
  doutReg = _RAND_41[63:0];
  _RAND_42 = {1{`RANDOM}};
  validReg = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  lruReg = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  wayReg = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  cacheEntryReg_valid = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  cacheEntryReg_tag = _RAND_46[26:0];
  _RAND_47 = {1{`RANDOM}};
  cacheEntryReg_line_words_0 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  cacheEntryReg_line_words_1 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  cacheEntryReg_line_words_2 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  cacheEntryReg_line_words_3 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  initCounter = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  burstCounter = _RAND_52[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BurstMemArbiter(
  input         clock,
  input         reset,
  input         io_in_0_wr,
  input  [31:0] io_in_0_addr,
  input  [63:0] io_in_0_din,
  output        io_in_0_burstDone,
  input         io_in_1_rd,
  input  [31:0] io_in_1_addr,
  output [63:0] io_in_1_dout,
  output        io_in_1_wait_n,
  output        io_in_1_valid,
  output        io_in_1_burstDone,
  input         io_in_2_wr,
  input  [31:0] io_in_2_addr,
  input  [7:0]  io_in_2_mask,
  input  [63:0] io_in_2_din,
  output        io_in_2_wait_n,
  input         io_in_3_rd,
  input         io_in_3_wr,
  input  [31:0] io_in_3_addr,
  input  [7:0]  io_in_3_mask,
  input  [63:0] io_in_3_din,
  output [63:0] io_in_3_dout,
  output        io_in_3_wait_n,
  output        io_in_3_valid,
  input  [7:0]  io_in_3_burstLength,
  output        io_in_3_burstDone,
  input         io_in_4_rd,
  input  [31:0] io_in_4_addr,
  output [63:0] io_in_4_dout,
  output        io_in_4_wait_n,
  output        io_in_4_valid,
  input  [7:0]  io_in_4_burstLength,
  output        io_in_4_burstDone,
  output        io_out_rd,
  output        io_out_wr,
  output [31:0] io_out_addr,
  output [7:0]  io_out_mask,
  output [63:0] io_out_din,
  input  [63:0] io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid,
  output [7:0]  io_out_burstLength,
  input         io_out_burstDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  busyReg; // @[BurstMemArbiter.scala 73:24]
  reg [4:0] indexReg; // @[BurstMemArbiter.scala 74:25]
  wire  _index_T_3 = io_in_3_rd | io_in_3_wr; // @[BurstMemArbiter.scala 77:65]
  wire [4:0] _index_enc_T = io_in_4_rd ? 5'h10 : 5'h0; // @[Mux.scala 47:70]
  wire [4:0] _index_enc_T_1 = _index_T_3 ? 5'h8 : _index_enc_T; // @[Mux.scala 47:70]
  wire [4:0] _index_enc_T_2 = io_in_2_wr ? 5'h4 : _index_enc_T_1; // @[Mux.scala 47:70]
  wire [4:0] _index_enc_T_3 = io_in_1_rd ? 5'h2 : _index_enc_T_2; // @[Mux.scala 47:70]
  wire [4:0] index_enc = io_in_0_wr ? 5'h1 : _index_enc_T_3; // @[Mux.scala 47:70]
  wire [4:0] index = {index_enc[4],index_enc[3],index_enc[2],index_enc[1],index_enc[0]}; // @[BurstMemArbiter.scala 77:78]
  wire [4:0] chosen = busyReg ? indexReg : index; // @[BurstMemArbiter.scala 80:19]
  wire  effectiveRequest = ~busyReg & (io_out_rd | io_out_wr) & io_out_wait_n; // @[BurstMemArbiter.scala 83:63]
  wire  _GEN_0 = effectiveRequest | busyReg; // @[BurstMemArbiter.scala 88:32 89:13 73:24]
  wire  io_out_anySelected = chosen[0] | chosen[1] | chosen[2] | chosen[3] | chosen[4]; // @[BurstMemIO.scala 316:45]
  wire [7:0] _io_out_mem_burstLength_T = chosen[0] ? 8'h1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_burstLength_T_1 = chosen[1] ? 8'h10 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_burstLength_T_2 = chosen[2] ? 8'h1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_burstLength_T_3 = chosen[3] ? io_in_3_burstLength : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_burstLength_T_4 = chosen[4] ? io_in_4_burstLength : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_burstLength_T_5 = _io_out_mem_burstLength_T | _io_out_mem_burstLength_T_1; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_burstLength_T_6 = _io_out_mem_burstLength_T_5 | _io_out_mem_burstLength_T_2; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_burstLength_T_7 = _io_out_mem_burstLength_T_6 | _io_out_mem_burstLength_T_3; // @[Mux.scala 27:73]
  wire [31:0] _io_out_mem_addr_T = chosen[0] ? io_in_0_addr : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_out_mem_addr_T_1 = chosen[1] ? io_in_1_addr : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_out_mem_addr_T_2 = chosen[2] ? io_in_2_addr : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_out_mem_addr_T_3 = chosen[3] ? io_in_3_addr : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_out_mem_addr_T_4 = chosen[4] ? io_in_4_addr : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_out_mem_addr_T_5 = _io_out_mem_addr_T | _io_out_mem_addr_T_1; // @[Mux.scala 27:73]
  wire [31:0] _io_out_mem_addr_T_6 = _io_out_mem_addr_T_5 | _io_out_mem_addr_T_2; // @[Mux.scala 27:73]
  wire [31:0] _io_out_mem_addr_T_7 = _io_out_mem_addr_T_6 | _io_out_mem_addr_T_3; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_mask_T = chosen[0] ? 8'hff : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_mask_T_2 = chosen[2] ? io_in_2_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_mask_T_3 = chosen[3] ? io_in_3_mask : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_mask_T_6 = _io_out_mem_mask_T | _io_out_mem_mask_T_2; // @[Mux.scala 27:73]
  wire [63:0] _io_out_mem_din_T = chosen[0] ? io_in_0_din : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_mem_din_T_2 = chosen[2] ? io_in_2_din : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_mem_din_T_3 = chosen[3] ? io_in_3_din : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_mem_din_T_6 = _io_out_mem_din_T | _io_out_mem_din_T_2; // @[Mux.scala 27:73]
  assign io_in_0_burstDone = chosen[0] & io_out_burstDone; // @[BurstMemIO.scala 327:34]
  assign io_in_1_dout = io_out_dout; // @[BurstMemIO.scala 317:19 BurstMemArbiter.scala 96:10]
  assign io_in_1_wait_n = (~io_out_anySelected | chosen[1]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_1_valid = chosen[1] & io_out_valid; // @[BurstMemIO.scala 326:30]
  assign io_in_1_burstDone = chosen[1] & io_out_burstDone; // @[BurstMemIO.scala 327:34]
  assign io_in_2_wait_n = (~io_out_anySelected | chosen[2]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_3_dout = io_out_dout; // @[BurstMemIO.scala 317:19 BurstMemArbiter.scala 96:10]
  assign io_in_3_wait_n = (~io_out_anySelected | chosen[3]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_3_valid = chosen[3] & io_out_valid; // @[BurstMemIO.scala 326:30]
  assign io_in_3_burstDone = chosen[3] & io_out_burstDone; // @[BurstMemIO.scala 327:34]
  assign io_in_4_dout = io_out_dout; // @[BurstMemIO.scala 317:19 BurstMemArbiter.scala 96:10]
  assign io_in_4_wait_n = (~io_out_anySelected | chosen[4]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_4_valid = chosen[4] & io_out_valid; // @[BurstMemIO.scala 326:30]
  assign io_in_4_burstDone = chosen[4] & io_out_burstDone; // @[BurstMemIO.scala 327:34]
  assign io_out_rd = chosen[1] & io_in_1_rd | chosen[3] & io_in_3_rd | chosen[4] & io_in_4_rd; // @[Mux.scala 27:73]
  assign io_out_wr = chosen[0] & io_in_0_wr | chosen[2] & io_in_2_wr | chosen[3] & io_in_3_wr; // @[Mux.scala 27:73]
  assign io_out_addr = _io_out_mem_addr_T_7 | _io_out_mem_addr_T_4; // @[Mux.scala 27:73]
  assign io_out_mask = _io_out_mem_mask_T_6 | _io_out_mem_mask_T_3; // @[Mux.scala 27:73]
  assign io_out_din = _io_out_mem_din_T_6 | _io_out_mem_din_T_3; // @[Mux.scala 27:73]
  assign io_out_burstLength = _io_out_mem_burstLength_T_7 | _io_out_mem_burstLength_T_4; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (reset) begin // @[BurstMemArbiter.scala 73:24]
      busyReg <= 1'h0; // @[BurstMemArbiter.scala 73:24]
    end else if (io_out_burstDone) begin // @[BurstMemArbiter.scala 86:26]
      busyReg <= 1'h0; // @[BurstMemArbiter.scala 87:13]
    end else begin
      busyReg <= _GEN_0;
    end
    if (reset) begin // @[BurstMemArbiter.scala 74:25]
      indexReg <= 5'h0; // @[BurstMemArbiter.scala 74:25]
    end else if (!(io_out_burstDone)) begin // @[BurstMemArbiter.scala 86:26]
      if (effectiveRequest) begin // @[BurstMemArbiter.scala 88:32]
        indexReg <= index; // @[BurstMemArbiter.scala 90:14]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busyReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  indexReg = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BurstMemArbiter_1(
  input         clock,
  input         reset,
  input         io_in_0_wr,
  input  [24:0] io_in_0_addr,
  input  [15:0] io_in_0_din,
  output        io_in_0_wait_n,
  output        io_in_0_burstDone,
  input         io_in_1_rd,
  input  [24:0] io_in_1_addr,
  output [15:0] io_in_1_dout,
  output        io_in_1_wait_n,
  output        io_in_1_valid,
  input         io_in_2_rd,
  input         io_in_2_wr,
  input  [24:0] io_in_2_addr,
  input  [15:0] io_in_2_din,
  output [15:0] io_in_2_dout,
  output        io_in_2_wait_n,
  output        io_in_2_valid,
  input         io_in_3_rd,
  input  [24:0] io_in_3_addr,
  output [15:0] io_in_3_dout,
  output        io_in_3_wait_n,
  output        io_in_3_valid,
  input         io_in_4_rd,
  input  [24:0] io_in_4_addr,
  output [15:0] io_in_4_dout,
  output        io_in_4_wait_n,
  output        io_in_4_valid,
  input         io_in_5_rd,
  input  [24:0] io_in_5_addr,
  output [15:0] io_in_5_dout,
  output        io_in_5_wait_n,
  output        io_in_5_valid,
  input         io_in_6_rd,
  input  [24:0] io_in_6_addr,
  output [15:0] io_in_6_dout,
  output        io_in_6_wait_n,
  output        io_in_6_valid,
  input         io_in_7_rd,
  input  [24:0] io_in_7_addr,
  output [15:0] io_in_7_dout,
  output        io_in_7_wait_n,
  output        io_in_7_valid,
  output        io_out_rd,
  output        io_out_wr,
  output [24:0] io_out_addr,
  output [15:0] io_out_din,
  input  [15:0] io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid,
  input         io_out_burstDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  busyReg; // @[BurstMemArbiter.scala 73:24]
  reg [7:0] indexReg; // @[BurstMemArbiter.scala 74:25]
  wire  _index_T_2 = io_in_2_rd | io_in_2_wr; // @[BurstMemArbiter.scala 77:65]
  wire [7:0] _index_enc_T = io_in_7_rd ? 8'h80 : 8'h0; // @[Mux.scala 47:70]
  wire [7:0] _index_enc_T_1 = io_in_6_rd ? 8'h40 : _index_enc_T; // @[Mux.scala 47:70]
  wire [7:0] _index_enc_T_2 = io_in_5_rd ? 8'h20 : _index_enc_T_1; // @[Mux.scala 47:70]
  wire [7:0] _index_enc_T_3 = io_in_4_rd ? 8'h10 : _index_enc_T_2; // @[Mux.scala 47:70]
  wire [7:0] _index_enc_T_4 = io_in_3_rd ? 8'h8 : _index_enc_T_3; // @[Mux.scala 47:70]
  wire [7:0] _index_enc_T_5 = _index_T_2 ? 8'h4 : _index_enc_T_4; // @[Mux.scala 47:70]
  wire [7:0] _index_enc_T_6 = io_in_1_rd ? 8'h2 : _index_enc_T_5; // @[Mux.scala 47:70]
  wire [7:0] index_enc = io_in_0_wr ? 8'h1 : _index_enc_T_6; // @[Mux.scala 47:70]
  wire [7:0] index = {index_enc[7],index_enc[6],index_enc[5],index_enc[4],index_enc[3],index_enc[2],index_enc[1],
    index_enc[0]}; // @[BurstMemArbiter.scala 77:78]
  wire [7:0] chosen = busyReg ? indexReg : index; // @[BurstMemArbiter.scala 80:19]
  wire  effectiveRequest = ~busyReg & (io_out_rd | io_out_wr) & io_out_wait_n; // @[BurstMemArbiter.scala 83:63]
  wire  _GEN_0 = effectiveRequest | busyReg; // @[BurstMemArbiter.scala 88:32 89:13 73:24]
  wire  io_out_anySelected = chosen[0] | chosen[1] | chosen[2] | chosen[3] | chosen[4] | chosen[5] | chosen[6] | chosen[
    7]; // @[BurstMemIO.scala 316:45]
  wire [24:0] _io_out_mem_addr_T = chosen[0] ? io_in_0_addr : 25'h0; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_1 = chosen[1] ? io_in_1_addr : 25'h0; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_2 = chosen[2] ? io_in_2_addr : 25'h0; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_3 = chosen[3] ? io_in_3_addr : 25'h0; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_4 = chosen[4] ? io_in_4_addr : 25'h0; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_5 = chosen[5] ? io_in_5_addr : 25'h0; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_6 = chosen[6] ? io_in_6_addr : 25'h0; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_7 = chosen[7] ? io_in_7_addr : 25'h0; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_8 = _io_out_mem_addr_T | _io_out_mem_addr_T_1; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_9 = _io_out_mem_addr_T_8 | _io_out_mem_addr_T_2; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_10 = _io_out_mem_addr_T_9 | _io_out_mem_addr_T_3; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_11 = _io_out_mem_addr_T_10 | _io_out_mem_addr_T_4; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_12 = _io_out_mem_addr_T_11 | _io_out_mem_addr_T_5; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_13 = _io_out_mem_addr_T_12 | _io_out_mem_addr_T_6; // @[Mux.scala 27:73]
  wire [15:0] _io_out_mem_din_T = chosen[0] ? io_in_0_din : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_out_mem_din_T_2 = chosen[2] ? io_in_2_din : 16'h0; // @[Mux.scala 27:73]
  assign io_in_0_wait_n = (~io_out_anySelected | chosen[0]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_0_burstDone = chosen[0] & io_out_burstDone; // @[BurstMemIO.scala 327:34]
  assign io_in_1_dout = io_out_dout; // @[BurstMemIO.scala 317:19 BurstMemArbiter.scala 96:10]
  assign io_in_1_wait_n = (~io_out_anySelected | chosen[1]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_1_valid = chosen[1] & io_out_valid; // @[BurstMemIO.scala 326:30]
  assign io_in_2_dout = io_out_dout; // @[BurstMemIO.scala 317:19 BurstMemArbiter.scala 96:10]
  assign io_in_2_wait_n = (~io_out_anySelected | chosen[2]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_2_valid = chosen[2] & io_out_valid; // @[BurstMemIO.scala 326:30]
  assign io_in_3_dout = io_out_dout; // @[BurstMemIO.scala 317:19 BurstMemArbiter.scala 96:10]
  assign io_in_3_wait_n = (~io_out_anySelected | chosen[3]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_3_valid = chosen[3] & io_out_valid; // @[BurstMemIO.scala 326:30]
  assign io_in_4_dout = io_out_dout; // @[BurstMemIO.scala 317:19 BurstMemArbiter.scala 96:10]
  assign io_in_4_wait_n = (~io_out_anySelected | chosen[4]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_4_valid = chosen[4] & io_out_valid; // @[BurstMemIO.scala 326:30]
  assign io_in_5_dout = io_out_dout; // @[BurstMemIO.scala 317:19 BurstMemArbiter.scala 96:10]
  assign io_in_5_wait_n = (~io_out_anySelected | chosen[5]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_5_valid = chosen[5] & io_out_valid; // @[BurstMemIO.scala 326:30]
  assign io_in_6_dout = io_out_dout; // @[BurstMemIO.scala 317:19 BurstMemArbiter.scala 96:10]
  assign io_in_6_wait_n = (~io_out_anySelected | chosen[6]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_6_valid = chosen[6] & io_out_valid; // @[BurstMemIO.scala 326:30]
  assign io_in_7_dout = io_out_dout; // @[BurstMemIO.scala 317:19 BurstMemArbiter.scala 96:10]
  assign io_in_7_wait_n = (~io_out_anySelected | chosen[7]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_7_valid = chosen[7] & io_out_valid; // @[BurstMemIO.scala 326:30]
  assign io_out_rd = chosen[1] & io_in_1_rd | chosen[2] & io_in_2_rd | chosen[3] & io_in_3_rd | chosen[4] & io_in_4_rd
     | chosen[5] & io_in_5_rd | chosen[6] & io_in_6_rd | chosen[7] & io_in_7_rd; // @[Mux.scala 27:73]
  assign io_out_wr = chosen[0] & io_in_0_wr | chosen[2] & io_in_2_wr; // @[Mux.scala 27:73]
  assign io_out_addr = _io_out_mem_addr_T_13 | _io_out_mem_addr_T_7; // @[Mux.scala 27:73]
  assign io_out_din = _io_out_mem_din_T | _io_out_mem_din_T_2; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (reset) begin // @[BurstMemArbiter.scala 73:24]
      busyReg <= 1'h0; // @[BurstMemArbiter.scala 73:24]
    end else if (io_out_burstDone) begin // @[BurstMemArbiter.scala 86:26]
      busyReg <= 1'h0; // @[BurstMemArbiter.scala 87:13]
    end else begin
      busyReg <= _GEN_0;
    end
    if (reset) begin // @[BurstMemArbiter.scala 74:25]
      indexReg <= 8'h0; // @[BurstMemArbiter.scala 74:25]
    end else if (!(io_out_burstDone)) begin // @[BurstMemArbiter.scala 86:26]
      if (effectiveRequest) begin // @[BurstMemArbiter.scala 88:32]
        indexReg <= index; // @[BurstMemArbiter.scala 90:14]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busyReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  indexReg = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncMemArbiter(
  input         clock,
  input         reset,
  input         io_in_0_rd,
  input         io_in_0_wr,
  input  [6:0]  io_in_0_addr,
  input  [15:0] io_in_0_din,
  output [15:0] io_in_0_dout,
  output        io_in_0_wait_n,
  output        io_in_0_valid,
  input         io_in_1_rd,
  input         io_in_1_wr,
  input  [6:0]  io_in_1_addr,
  input  [15:0] io_in_1_din,
  output [15:0] io_in_1_dout,
  output        io_in_1_wait_n,
  output        io_in_1_valid,
  output        io_out_rd,
  output        io_out_wr,
  output [6:0]  io_out_addr,
  output [15:0] io_out_din,
  input  [15:0] io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  busyReg; // @[AsyncMemArbiter.scala 73:24]
  reg [1:0] indexReg; // @[AsyncMemArbiter.scala 74:25]
  wire  _index_T = io_in_0_rd | io_in_0_wr; // @[AsyncMemArbiter.scala 77:65]
  wire  _index_T_1 = io_in_1_rd | io_in_1_wr; // @[AsyncMemArbiter.scala 77:65]
  wire [1:0] _index_enc_T = _index_T_1 ? 2'h2 : 2'h0; // @[Mux.scala 47:70]
  wire [1:0] index_enc = _index_T ? 2'h1 : _index_enc_T; // @[Mux.scala 47:70]
  wire [1:0] index = {index_enc[1],index_enc[0]}; // @[AsyncMemArbiter.scala 77:78]
  wire [1:0] chosen = busyReg ? indexReg : index; // @[AsyncMemArbiter.scala 80:19]
  wire  effectiveRequest = ~busyReg & io_out_rd & io_out_wait_n; // @[AsyncMemArbiter.scala 83:48]
  wire  _GEN_0 = effectiveRequest | busyReg; // @[AsyncMemArbiter.scala 88:32 89:13 73:24]
  wire  io_out_anySelected = chosen[0] | chosen[1]; // @[AsyncMemIO.scala 354:45]
  wire [6:0] _io_out_mem_addr_T = chosen[0] ? io_in_0_addr : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_out_mem_addr_T_1 = chosen[1] ? io_in_1_addr : 7'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_out_mem_din_T = chosen[0] ? io_in_0_din : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_out_mem_din_T_1 = chosen[1] ? io_in_1_din : 16'h0; // @[Mux.scala 27:73]
  assign io_in_0_dout = io_out_dout; // @[AsyncMemIO.scala 355:19 AsyncMemArbiter.scala 96:10]
  assign io_in_0_wait_n = (~io_out_anySelected | chosen[0]) & io_out_wait_n; // @[AsyncMemIO.scala 362:49]
  assign io_in_0_valid = chosen[0] & io_out_valid; // @[AsyncMemIO.scala 363:30]
  assign io_in_1_dout = io_out_dout; // @[AsyncMemIO.scala 355:19 AsyncMemArbiter.scala 96:10]
  assign io_in_1_wait_n = (~io_out_anySelected | chosen[1]) & io_out_wait_n; // @[AsyncMemIO.scala 362:49]
  assign io_in_1_valid = chosen[1] & io_out_valid; // @[AsyncMemIO.scala 363:30]
  assign io_out_rd = chosen[0] & io_in_0_rd | chosen[1] & io_in_1_rd; // @[Mux.scala 27:73]
  assign io_out_wr = chosen[0] & io_in_0_wr | chosen[1] & io_in_1_wr; // @[Mux.scala 27:73]
  assign io_out_addr = _io_out_mem_addr_T | _io_out_mem_addr_T_1; // @[Mux.scala 27:73]
  assign io_out_din = _io_out_mem_din_T | _io_out_mem_din_T_1; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (reset) begin // @[AsyncMemArbiter.scala 73:24]
      busyReg <= 1'h0; // @[AsyncMemArbiter.scala 73:24]
    end else if (io_out_valid) begin // @[AsyncMemArbiter.scala 86:22]
      busyReg <= 1'h0; // @[AsyncMemArbiter.scala 87:13]
    end else begin
      busyReg <= _GEN_0;
    end
    if (reset) begin // @[AsyncMemArbiter.scala 74:25]
      indexReg <= 2'h0; // @[AsyncMemArbiter.scala 74:25]
    end else if (!(io_out_valid)) begin // @[AsyncMemArbiter.scala 86:22]
      if (effectiveRequest) begin // @[AsyncMemArbiter.scala 88:32]
        indexReg <= index; // @[AsyncMemArbiter.scala 90:14]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busyReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  indexReg = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemSys(
  input         clock,
  input         reset,
  input  [31:0] io_gameConfig_eepromOffset,
  input  [31:0] io_gameConfig_sound_0_romOffset,
  input  [31:0] io_gameConfig_sound_1_romOffset,
  input  [31:0] io_gameConfig_layer_0_romOffset,
  input  [31:0] io_gameConfig_layer_1_romOffset,
  input  [31:0] io_gameConfig_layer_2_romOffset,
  input  [31:0] io_gameConfig_sprite_romOffset,
  input         io_prog_rom_wr,
  input  [26:0] io_prog_rom_addr,
  input  [15:0] io_prog_rom_din,
  output        io_prog_rom_wait_n,
  input         io_prog_nvram_rd,
  input         io_prog_nvram_wr,
  input  [26:0] io_prog_nvram_addr,
  input  [15:0] io_prog_nvram_din,
  output [15:0] io_prog_nvram_dout,
  output        io_prog_nvram_wait_n,
  output        io_prog_nvram_valid,
  input         io_prog_done,
  input         io_progRom_rd,
  input  [19:0] io_progRom_addr,
  output [15:0] io_progRom_dout,
  output        io_progRom_wait_n,
  output        io_progRom_valid,
  input         io_eeprom_rd,
  input         io_eeprom_wr,
  input  [6:0]  io_eeprom_addr,
  input  [15:0] io_eeprom_din,
  output [15:0] io_eeprom_dout,
  output        io_eeprom_wait_n,
  output        io_eeprom_valid,
  input         io_soundRom_0_rd,
  input  [24:0] io_soundRom_0_addr,
  output [7:0]  io_soundRom_0_dout,
  output        io_soundRom_0_wait_n,
  output        io_soundRom_0_valid,
  input         io_soundRom_1_rd,
  input  [24:0] io_soundRom_1_addr,
  output [7:0]  io_soundRom_1_dout,
  output        io_soundRom_1_wait_n,
  output        io_soundRom_1_valid,
  input         io_layerTileRom_0_rd,
  input  [31:0] io_layerTileRom_0_addr,
  output [63:0] io_layerTileRom_0_dout,
  output        io_layerTileRom_0_wait_n,
  output        io_layerTileRom_0_valid,
  input         io_layerTileRom_1_rd,
  input  [31:0] io_layerTileRom_1_addr,
  output [63:0] io_layerTileRom_1_dout,
  output        io_layerTileRom_1_wait_n,
  output        io_layerTileRom_1_valid,
  input         io_layerTileRom_2_rd,
  input  [31:0] io_layerTileRom_2_addr,
  output [63:0] io_layerTileRom_2_dout,
  output        io_layerTileRom_2_wait_n,
  output        io_layerTileRom_2_valid,
  input         io_spriteTileRom_rd,
  input  [31:0] io_spriteTileRom_addr,
  output [63:0] io_spriteTileRom_dout,
  output        io_spriteTileRom_wait_n,
  output        io_spriteTileRom_valid,
  input  [7:0]  io_spriteTileRom_burstLength,
  output        io_spriteTileRom_burstDone,
  output        io_ddr_rd,
  output        io_ddr_wr,
  output [31:0] io_ddr_addr,
  output [7:0]  io_ddr_mask,
  output [63:0] io_ddr_din,
  input  [63:0] io_ddr_dout,
  input         io_ddr_wait_n,
  input         io_ddr_valid,
  output [7:0]  io_ddr_burstLength,
  input         io_ddr_burstDone,
  output        io_sdram_rd,
  output        io_sdram_wr,
  output [24:0] io_sdram_addr,
  output [15:0] io_sdram_din,
  input  [15:0] io_sdram_dout,
  input         io_sdram_wait_n,
  input         io_sdram_valid,
  input         io_sdram_burstDone,
  input         io_spriteFrameBuffer_rd,
  input         io_spriteFrameBuffer_wr,
  input  [31:0] io_spriteFrameBuffer_addr,
  input  [7:0]  io_spriteFrameBuffer_mask,
  input  [63:0] io_spriteFrameBuffer_din,
  output [63:0] io_spriteFrameBuffer_dout,
  output        io_spriteFrameBuffer_wait_n,
  output        io_spriteFrameBuffer_valid,
  input  [7:0]  io_spriteFrameBuffer_burstLength,
  output        io_spriteFrameBuffer_burstDone,
  input         io_systemFrameBuffer_wr,
  input  [31:0] io_systemFrameBuffer_addr,
  input  [7:0]  io_systemFrameBuffer_mask,
  input  [63:0] io_systemFrameBuffer_din,
  output        io_systemFrameBuffer_wait_n,
  output        io_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  ddrDownloadBuffer_clock; // @[MemSys.scala 82:33]
  wire  ddrDownloadBuffer_reset; // @[MemSys.scala 82:33]
  wire  ddrDownloadBuffer_io_in_wr; // @[MemSys.scala 82:33]
  wire [26:0] ddrDownloadBuffer_io_in_addr; // @[MemSys.scala 82:33]
  wire [15:0] ddrDownloadBuffer_io_in_din; // @[MemSys.scala 82:33]
  wire  ddrDownloadBuffer_io_out_wr; // @[MemSys.scala 82:33]
  wire [31:0] ddrDownloadBuffer_io_out_addr; // @[MemSys.scala 82:33]
  wire [63:0] ddrDownloadBuffer_io_out_din; // @[MemSys.scala 82:33]
  wire  ddrDownloadBuffer_io_out_burstDone; // @[MemSys.scala 82:33]
  wire  sdramDownloadBuffer_clock; // @[MemSys.scala 92:35]
  wire  sdramDownloadBuffer_reset; // @[MemSys.scala 92:35]
  wire  sdramDownloadBuffer_io_in_wr; // @[MemSys.scala 92:35]
  wire [31:0] sdramDownloadBuffer_io_in_addr; // @[MemSys.scala 92:35]
  wire [63:0] sdramDownloadBuffer_io_in_din; // @[MemSys.scala 92:35]
  wire  sdramDownloadBuffer_io_in_wait_n; // @[MemSys.scala 92:35]
  wire  sdramDownloadBuffer_io_out_wr; // @[MemSys.scala 92:35]
  wire [24:0] sdramDownloadBuffer_io_out_addr; // @[MemSys.scala 92:35]
  wire [15:0] sdramDownloadBuffer_io_out_din; // @[MemSys.scala 92:35]
  wire  sdramDownloadBuffer_io_out_wait_n; // @[MemSys.scala 92:35]
  wire  sdramDownloadBuffer_io_out_burstDone; // @[MemSys.scala 92:35]
  wire  copyDma_clock; // @[MemSys.scala 102:23]
  wire  copyDma_reset; // @[MemSys.scala 102:23]
  wire  copyDma_io_start; // @[MemSys.scala 102:23]
  wire  copyDma_io_busy; // @[MemSys.scala 102:23]
  wire  copyDma_io_in_rd; // @[MemSys.scala 102:23]
  wire [31:0] copyDma_io_in_addr; // @[MemSys.scala 102:23]
  wire [63:0] copyDma_io_in_dout; // @[MemSys.scala 102:23]
  wire  copyDma_io_in_wait_n; // @[MemSys.scala 102:23]
  wire  copyDma_io_in_valid; // @[MemSys.scala 102:23]
  wire  copyDma_io_in_burstDone; // @[MemSys.scala 102:23]
  wire  copyDma_io_out_wr; // @[MemSys.scala 102:23]
  wire [31:0] copyDma_io_out_addr; // @[MemSys.scala 102:23]
  wire [63:0] copyDma_io_out_din; // @[MemSys.scala 102:23]
  wire  copyDma_io_out_wait_n; // @[MemSys.scala 102:23]
  wire  progRomCache_clock; // @[MemSys.scala 107:28]
  wire  progRomCache_reset; // @[MemSys.scala 107:28]
  wire  progRomCache_io_enable; // @[MemSys.scala 107:28]
  wire  progRomCache_io_in_rd; // @[MemSys.scala 107:28]
  wire [19:0] progRomCache_io_in_addr; // @[MemSys.scala 107:28]
  wire [15:0] progRomCache_io_in_dout; // @[MemSys.scala 107:28]
  wire  progRomCache_io_in_wait_n; // @[MemSys.scala 107:28]
  wire  progRomCache_io_in_valid; // @[MemSys.scala 107:28]
  wire  progRomCache_io_out_rd; // @[MemSys.scala 107:28]
  wire [24:0] progRomCache_io_out_addr; // @[MemSys.scala 107:28]
  wire [15:0] progRomCache_io_out_dout; // @[MemSys.scala 107:28]
  wire  progRomCache_io_out_wait_n; // @[MemSys.scala 107:28]
  wire  progRomCache_io_out_valid; // @[MemSys.scala 107:28]
  wire  eepromCache_clock; // @[MemSys.scala 120:27]
  wire  eepromCache_reset; // @[MemSys.scala 120:27]
  wire  eepromCache_io_enable; // @[MemSys.scala 120:27]
  wire  eepromCache_io_in_rd; // @[MemSys.scala 120:27]
  wire  eepromCache_io_in_wr; // @[MemSys.scala 120:27]
  wire [6:0] eepromCache_io_in_addr; // @[MemSys.scala 120:27]
  wire [15:0] eepromCache_io_in_din; // @[MemSys.scala 120:27]
  wire [15:0] eepromCache_io_in_dout; // @[MemSys.scala 120:27]
  wire  eepromCache_io_in_wait_n; // @[MemSys.scala 120:27]
  wire  eepromCache_io_in_valid; // @[MemSys.scala 120:27]
  wire  eepromCache_io_out_rd; // @[MemSys.scala 120:27]
  wire  eepromCache_io_out_wr; // @[MemSys.scala 120:27]
  wire [24:0] eepromCache_io_out_addr; // @[MemSys.scala 120:27]
  wire [15:0] eepromCache_io_out_din; // @[MemSys.scala 120:27]
  wire [15:0] eepromCache_io_out_dout; // @[MemSys.scala 120:27]
  wire  eepromCache_io_out_wait_n; // @[MemSys.scala 120:27]
  wire  eepromCache_io_out_valid; // @[MemSys.scala 120:27]
  wire  soundRomCache_0_clock; // @[MemSys.scala 133:19]
  wire  soundRomCache_0_reset; // @[MemSys.scala 133:19]
  wire  soundRomCache_0_io_enable; // @[MemSys.scala 133:19]
  wire  soundRomCache_0_io_in_rd; // @[MemSys.scala 133:19]
  wire [24:0] soundRomCache_0_io_in_addr; // @[MemSys.scala 133:19]
  wire [7:0] soundRomCache_0_io_in_dout; // @[MemSys.scala 133:19]
  wire  soundRomCache_0_io_in_wait_n; // @[MemSys.scala 133:19]
  wire  soundRomCache_0_io_in_valid; // @[MemSys.scala 133:19]
  wire  soundRomCache_0_io_out_rd; // @[MemSys.scala 133:19]
  wire [24:0] soundRomCache_0_io_out_addr; // @[MemSys.scala 133:19]
  wire [15:0] soundRomCache_0_io_out_dout; // @[MemSys.scala 133:19]
  wire  soundRomCache_0_io_out_wait_n; // @[MemSys.scala 133:19]
  wire  soundRomCache_0_io_out_valid; // @[MemSys.scala 133:19]
  wire  soundRomCache_1_clock; // @[MemSys.scala 133:19]
  wire  soundRomCache_1_reset; // @[MemSys.scala 133:19]
  wire  soundRomCache_1_io_enable; // @[MemSys.scala 133:19]
  wire  soundRomCache_1_io_in_rd; // @[MemSys.scala 133:19]
  wire [24:0] soundRomCache_1_io_in_addr; // @[MemSys.scala 133:19]
  wire [7:0] soundRomCache_1_io_in_dout; // @[MemSys.scala 133:19]
  wire  soundRomCache_1_io_in_wait_n; // @[MemSys.scala 133:19]
  wire  soundRomCache_1_io_in_valid; // @[MemSys.scala 133:19]
  wire  soundRomCache_1_io_out_rd; // @[MemSys.scala 133:19]
  wire [24:0] soundRomCache_1_io_out_addr; // @[MemSys.scala 133:19]
  wire [15:0] soundRomCache_1_io_out_dout; // @[MemSys.scala 133:19]
  wire  soundRomCache_1_io_out_wait_n; // @[MemSys.scala 133:19]
  wire  soundRomCache_1_io_out_valid; // @[MemSys.scala 133:19]
  wire  layerRomCache_0_clock; // @[MemSys.scala 149:19]
  wire  layerRomCache_0_reset; // @[MemSys.scala 149:19]
  wire  layerRomCache_0_io_enable; // @[MemSys.scala 149:19]
  wire  layerRomCache_0_io_in_rd; // @[MemSys.scala 149:19]
  wire [31:0] layerRomCache_0_io_in_addr; // @[MemSys.scala 149:19]
  wire [63:0] layerRomCache_0_io_in_dout; // @[MemSys.scala 149:19]
  wire  layerRomCache_0_io_in_wait_n; // @[MemSys.scala 149:19]
  wire  layerRomCache_0_io_in_valid; // @[MemSys.scala 149:19]
  wire  layerRomCache_0_io_out_rd; // @[MemSys.scala 149:19]
  wire [24:0] layerRomCache_0_io_out_addr; // @[MemSys.scala 149:19]
  wire [15:0] layerRomCache_0_io_out_dout; // @[MemSys.scala 149:19]
  wire  layerRomCache_0_io_out_wait_n; // @[MemSys.scala 149:19]
  wire  layerRomCache_0_io_out_valid; // @[MemSys.scala 149:19]
  wire  layerRomCache_1_clock; // @[MemSys.scala 149:19]
  wire  layerRomCache_1_reset; // @[MemSys.scala 149:19]
  wire  layerRomCache_1_io_enable; // @[MemSys.scala 149:19]
  wire  layerRomCache_1_io_in_rd; // @[MemSys.scala 149:19]
  wire [31:0] layerRomCache_1_io_in_addr; // @[MemSys.scala 149:19]
  wire [63:0] layerRomCache_1_io_in_dout; // @[MemSys.scala 149:19]
  wire  layerRomCache_1_io_in_wait_n; // @[MemSys.scala 149:19]
  wire  layerRomCache_1_io_in_valid; // @[MemSys.scala 149:19]
  wire  layerRomCache_1_io_out_rd; // @[MemSys.scala 149:19]
  wire [24:0] layerRomCache_1_io_out_addr; // @[MemSys.scala 149:19]
  wire [15:0] layerRomCache_1_io_out_dout; // @[MemSys.scala 149:19]
  wire  layerRomCache_1_io_out_wait_n; // @[MemSys.scala 149:19]
  wire  layerRomCache_1_io_out_valid; // @[MemSys.scala 149:19]
  wire  layerRomCache_2_clock; // @[MemSys.scala 149:19]
  wire  layerRomCache_2_reset; // @[MemSys.scala 149:19]
  wire  layerRomCache_2_io_enable; // @[MemSys.scala 149:19]
  wire  layerRomCache_2_io_in_rd; // @[MemSys.scala 149:19]
  wire [31:0] layerRomCache_2_io_in_addr; // @[MemSys.scala 149:19]
  wire [63:0] layerRomCache_2_io_in_dout; // @[MemSys.scala 149:19]
  wire  layerRomCache_2_io_in_wait_n; // @[MemSys.scala 149:19]
  wire  layerRomCache_2_io_in_valid; // @[MemSys.scala 149:19]
  wire  layerRomCache_2_io_out_rd; // @[MemSys.scala 149:19]
  wire [24:0] layerRomCache_2_io_out_addr; // @[MemSys.scala 149:19]
  wire [15:0] layerRomCache_2_io_out_dout; // @[MemSys.scala 149:19]
  wire  layerRomCache_2_io_out_wait_n; // @[MemSys.scala 149:19]
  wire  layerRomCache_2_io_out_valid; // @[MemSys.scala 149:19]
  wire  ddrArbiter_clock; // @[MemSys.scala 164:26]
  wire  ddrArbiter_reset; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_0_wr; // @[MemSys.scala 164:26]
  wire [31:0] ddrArbiter_io_in_0_addr; // @[MemSys.scala 164:26]
  wire [63:0] ddrArbiter_io_in_0_din; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_0_burstDone; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_1_rd; // @[MemSys.scala 164:26]
  wire [31:0] ddrArbiter_io_in_1_addr; // @[MemSys.scala 164:26]
  wire [63:0] ddrArbiter_io_in_1_dout; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_1_wait_n; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_1_valid; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_1_burstDone; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_2_wr; // @[MemSys.scala 164:26]
  wire [31:0] ddrArbiter_io_in_2_addr; // @[MemSys.scala 164:26]
  wire [7:0] ddrArbiter_io_in_2_mask; // @[MemSys.scala 164:26]
  wire [63:0] ddrArbiter_io_in_2_din; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_2_wait_n; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_3_rd; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_3_wr; // @[MemSys.scala 164:26]
  wire [31:0] ddrArbiter_io_in_3_addr; // @[MemSys.scala 164:26]
  wire [7:0] ddrArbiter_io_in_3_mask; // @[MemSys.scala 164:26]
  wire [63:0] ddrArbiter_io_in_3_din; // @[MemSys.scala 164:26]
  wire [63:0] ddrArbiter_io_in_3_dout; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_3_wait_n; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_3_valid; // @[MemSys.scala 164:26]
  wire [7:0] ddrArbiter_io_in_3_burstLength; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_3_burstDone; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_4_rd; // @[MemSys.scala 164:26]
  wire [31:0] ddrArbiter_io_in_4_addr; // @[MemSys.scala 164:26]
  wire [63:0] ddrArbiter_io_in_4_dout; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_4_wait_n; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_4_valid; // @[MemSys.scala 164:26]
  wire [7:0] ddrArbiter_io_in_4_burstLength; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_in_4_burstDone; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_out_rd; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_out_wr; // @[MemSys.scala 164:26]
  wire [31:0] ddrArbiter_io_out_addr; // @[MemSys.scala 164:26]
  wire [7:0] ddrArbiter_io_out_mask; // @[MemSys.scala 164:26]
  wire [63:0] ddrArbiter_io_out_din; // @[MemSys.scala 164:26]
  wire [63:0] ddrArbiter_io_out_dout; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_out_wait_n; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_out_valid; // @[MemSys.scala 164:26]
  wire [7:0] ddrArbiter_io_out_burstLength; // @[MemSys.scala 164:26]
  wire  ddrArbiter_io_out_burstDone; // @[MemSys.scala 164:26]
  wire  sdramArbiter_clock; // @[MemSys.scala 174:28]
  wire  sdramArbiter_reset; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_0_wr; // @[MemSys.scala 174:28]
  wire [24:0] sdramArbiter_io_in_0_addr; // @[MemSys.scala 174:28]
  wire [15:0] sdramArbiter_io_in_0_din; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_0_wait_n; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_0_burstDone; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_1_rd; // @[MemSys.scala 174:28]
  wire [24:0] sdramArbiter_io_in_1_addr; // @[MemSys.scala 174:28]
  wire [15:0] sdramArbiter_io_in_1_dout; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_1_wait_n; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_1_valid; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_2_rd; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_2_wr; // @[MemSys.scala 174:28]
  wire [24:0] sdramArbiter_io_in_2_addr; // @[MemSys.scala 174:28]
  wire [15:0] sdramArbiter_io_in_2_din; // @[MemSys.scala 174:28]
  wire [15:0] sdramArbiter_io_in_2_dout; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_2_wait_n; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_2_valid; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_3_rd; // @[MemSys.scala 174:28]
  wire [24:0] sdramArbiter_io_in_3_addr; // @[MemSys.scala 174:28]
  wire [15:0] sdramArbiter_io_in_3_dout; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_3_wait_n; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_3_valid; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_4_rd; // @[MemSys.scala 174:28]
  wire [24:0] sdramArbiter_io_in_4_addr; // @[MemSys.scala 174:28]
  wire [15:0] sdramArbiter_io_in_4_dout; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_4_wait_n; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_4_valid; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_5_rd; // @[MemSys.scala 174:28]
  wire [24:0] sdramArbiter_io_in_5_addr; // @[MemSys.scala 174:28]
  wire [15:0] sdramArbiter_io_in_5_dout; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_5_wait_n; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_5_valid; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_6_rd; // @[MemSys.scala 174:28]
  wire [24:0] sdramArbiter_io_in_6_addr; // @[MemSys.scala 174:28]
  wire [15:0] sdramArbiter_io_in_6_dout; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_6_wait_n; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_6_valid; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_7_rd; // @[MemSys.scala 174:28]
  wire [24:0] sdramArbiter_io_in_7_addr; // @[MemSys.scala 174:28]
  wire [15:0] sdramArbiter_io_in_7_dout; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_7_wait_n; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_in_7_valid; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_out_rd; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_out_wr; // @[MemSys.scala 174:28]
  wire [24:0] sdramArbiter_io_out_addr; // @[MemSys.scala 174:28]
  wire [15:0] sdramArbiter_io_out_din; // @[MemSys.scala 174:28]
  wire [15:0] sdramArbiter_io_out_dout; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_out_wait_n; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_out_valid; // @[MemSys.scala 174:28]
  wire  sdramArbiter_io_out_burstDone; // @[MemSys.scala 174:28]
  wire  nvramArbiter_clock; // @[MemSys.scala 187:28]
  wire  nvramArbiter_reset; // @[MemSys.scala 187:28]
  wire  nvramArbiter_io_in_0_rd; // @[MemSys.scala 187:28]
  wire  nvramArbiter_io_in_0_wr; // @[MemSys.scala 187:28]
  wire [6:0] nvramArbiter_io_in_0_addr; // @[MemSys.scala 187:28]
  wire [15:0] nvramArbiter_io_in_0_din; // @[MemSys.scala 187:28]
  wire [15:0] nvramArbiter_io_in_0_dout; // @[MemSys.scala 187:28]
  wire  nvramArbiter_io_in_0_wait_n; // @[MemSys.scala 187:28]
  wire  nvramArbiter_io_in_0_valid; // @[MemSys.scala 187:28]
  wire  nvramArbiter_io_in_1_rd; // @[MemSys.scala 187:28]
  wire  nvramArbiter_io_in_1_wr; // @[MemSys.scala 187:28]
  wire [6:0] nvramArbiter_io_in_1_addr; // @[MemSys.scala 187:28]
  wire [15:0] nvramArbiter_io_in_1_din; // @[MemSys.scala 187:28]
  wire [15:0] nvramArbiter_io_in_1_dout; // @[MemSys.scala 187:28]
  wire  nvramArbiter_io_in_1_wait_n; // @[MemSys.scala 187:28]
  wire  nvramArbiter_io_in_1_valid; // @[MemSys.scala 187:28]
  wire  nvramArbiter_io_out_rd; // @[MemSys.scala 187:28]
  wire  nvramArbiter_io_out_wr; // @[MemSys.scala 187:28]
  wire [6:0] nvramArbiter_io_out_addr; // @[MemSys.scala 187:28]
  wire [15:0] nvramArbiter_io_out_din; // @[MemSys.scala 187:28]
  wire [15:0] nvramArbiter_io_out_dout; // @[MemSys.scala 187:28]
  wire  nvramArbiter_io_out_wait_n; // @[MemSys.scala 187:28]
  wire  nvramArbiter_io_out_valid; // @[MemSys.scala 187:28]
  wire [31:0] _mem_T_5 = io_spriteTileRom_addr + io_gameConfig_sprite_romOffset; // @[MemSys.scala 170:32]
  wire [31:0] _GEN_2 = {{7'd0}, progRomCache_io_out_addr}; // @[MemSys.scala 177:35]
  wire [32:0] _mem_T_8 = {{1'd0}, _GEN_2}; // @[MemSys.scala 177:35]
  wire [31:0] _GEN_4 = {{7'd0}, eepromCache_io_out_addr}; // @[MemSys.scala 178:34]
  wire [31:0] _mem_T_11 = _GEN_4 + io_gameConfig_eepromOffset; // @[MemSys.scala 178:34]
  wire [31:0] _GEN_6 = {{7'd0}, soundRomCache_0_io_out_addr}; // @[MemSys.scala 179:39]
  wire [31:0] _mem_T_13 = _GEN_6 + io_gameConfig_sound_0_romOffset; // @[MemSys.scala 179:39]
  wire [31:0] _GEN_8 = {{7'd0}, soundRomCache_1_io_out_addr}; // @[MemSys.scala 180:39]
  wire [31:0] _mem_T_15 = _GEN_8 + io_gameConfig_sound_1_romOffset; // @[MemSys.scala 180:39]
  wire [31:0] _GEN_10 = {{7'd0}, layerRomCache_0_io_out_addr}; // @[MemSys.scala 181:39]
  wire [31:0] _mem_T_17 = _GEN_10 + io_gameConfig_layer_0_romOffset; // @[MemSys.scala 181:39]
  wire [31:0] _GEN_12 = {{7'd0}, layerRomCache_1_io_out_addr}; // @[MemSys.scala 182:39]
  wire [31:0] _mem_T_19 = _GEN_12 + io_gameConfig_layer_1_romOffset; // @[MemSys.scala 182:39]
  wire [31:0] _GEN_14 = {{7'd0}, layerRomCache_2_io_out_addr}; // @[MemSys.scala 183:39]
  wire [31:0] _mem_T_21 = _GEN_14 + io_gameConfig_layer_2_romOffset; // @[MemSys.scala 183:39]
  reg  io_ready_REG; // @[Util.scala 165:45]
  wire  _io_ready_T_1 = ~copyDma_io_busy & io_ready_REG; // @[Util.scala 165:35]
  reg  io_ready_enableReg; // @[Util.scala 218:28]
  wire  _GEN_0 = _io_ready_T_1 | io_ready_enableReg; // @[Util.scala 218:28 219:{54,66}]
  BurstBuffer ddrDownloadBuffer ( // @[MemSys.scala 82:33]
    .clock(ddrDownloadBuffer_clock),
    .reset(ddrDownloadBuffer_reset),
    .io_in_wr(ddrDownloadBuffer_io_in_wr),
    .io_in_addr(ddrDownloadBuffer_io_in_addr),
    .io_in_din(ddrDownloadBuffer_io_in_din),
    .io_out_wr(ddrDownloadBuffer_io_out_wr),
    .io_out_addr(ddrDownloadBuffer_io_out_addr),
    .io_out_din(ddrDownloadBuffer_io_out_din),
    .io_out_burstDone(ddrDownloadBuffer_io_out_burstDone)
  );
  BurstBuffer_1 sdramDownloadBuffer ( // @[MemSys.scala 92:35]
    .clock(sdramDownloadBuffer_clock),
    .reset(sdramDownloadBuffer_reset),
    .io_in_wr(sdramDownloadBuffer_io_in_wr),
    .io_in_addr(sdramDownloadBuffer_io_in_addr),
    .io_in_din(sdramDownloadBuffer_io_in_din),
    .io_in_wait_n(sdramDownloadBuffer_io_in_wait_n),
    .io_out_wr(sdramDownloadBuffer_io_out_wr),
    .io_out_addr(sdramDownloadBuffer_io_out_addr),
    .io_out_din(sdramDownloadBuffer_io_out_din),
    .io_out_wait_n(sdramDownloadBuffer_io_out_wait_n),
    .io_out_burstDone(sdramDownloadBuffer_io_out_burstDone)
  );
  BurstReadDMA copyDma ( // @[MemSys.scala 102:23]
    .clock(copyDma_clock),
    .reset(copyDma_reset),
    .io_start(copyDma_io_start),
    .io_busy(copyDma_io_busy),
    .io_in_rd(copyDma_io_in_rd),
    .io_in_addr(copyDma_io_in_addr),
    .io_in_dout(copyDma_io_in_dout),
    .io_in_wait_n(copyDma_io_in_wait_n),
    .io_in_valid(copyDma_io_in_valid),
    .io_in_burstDone(copyDma_io_in_burstDone),
    .io_out_wr(copyDma_io_out_wr),
    .io_out_addr(copyDma_io_out_addr),
    .io_out_din(copyDma_io_out_din),
    .io_out_wait_n(copyDma_io_out_wait_n)
  );
  ReadCache progRomCache ( // @[MemSys.scala 107:28]
    .clock(progRomCache_clock),
    .reset(progRomCache_reset),
    .io_enable(progRomCache_io_enable),
    .io_in_rd(progRomCache_io_in_rd),
    .io_in_addr(progRomCache_io_in_addr),
    .io_in_dout(progRomCache_io_in_dout),
    .io_in_wait_n(progRomCache_io_in_wait_n),
    .io_in_valid(progRomCache_io_in_valid),
    .io_out_rd(progRomCache_io_out_rd),
    .io_out_addr(progRomCache_io_out_addr),
    .io_out_dout(progRomCache_io_out_dout),
    .io_out_wait_n(progRomCache_io_out_wait_n),
    .io_out_valid(progRomCache_io_out_valid)
  );
  Cache eepromCache ( // @[MemSys.scala 120:27]
    .clock(eepromCache_clock),
    .reset(eepromCache_reset),
    .io_enable(eepromCache_io_enable),
    .io_in_rd(eepromCache_io_in_rd),
    .io_in_wr(eepromCache_io_in_wr),
    .io_in_addr(eepromCache_io_in_addr),
    .io_in_din(eepromCache_io_in_din),
    .io_in_dout(eepromCache_io_in_dout),
    .io_in_wait_n(eepromCache_io_in_wait_n),
    .io_in_valid(eepromCache_io_in_valid),
    .io_out_rd(eepromCache_io_out_rd),
    .io_out_wr(eepromCache_io_out_wr),
    .io_out_addr(eepromCache_io_out_addr),
    .io_out_din(eepromCache_io_out_din),
    .io_out_dout(eepromCache_io_out_dout),
    .io_out_wait_n(eepromCache_io_out_wait_n),
    .io_out_valid(eepromCache_io_out_valid)
  );
  ReadCache_1 soundRomCache_0 ( // @[MemSys.scala 133:19]
    .clock(soundRomCache_0_clock),
    .reset(soundRomCache_0_reset),
    .io_enable(soundRomCache_0_io_enable),
    .io_in_rd(soundRomCache_0_io_in_rd),
    .io_in_addr(soundRomCache_0_io_in_addr),
    .io_in_dout(soundRomCache_0_io_in_dout),
    .io_in_wait_n(soundRomCache_0_io_in_wait_n),
    .io_in_valid(soundRomCache_0_io_in_valid),
    .io_out_rd(soundRomCache_0_io_out_rd),
    .io_out_addr(soundRomCache_0_io_out_addr),
    .io_out_dout(soundRomCache_0_io_out_dout),
    .io_out_wait_n(soundRomCache_0_io_out_wait_n),
    .io_out_valid(soundRomCache_0_io_out_valid)
  );
  ReadCache_1 soundRomCache_1 ( // @[MemSys.scala 133:19]
    .clock(soundRomCache_1_clock),
    .reset(soundRomCache_1_reset),
    .io_enable(soundRomCache_1_io_enable),
    .io_in_rd(soundRomCache_1_io_in_rd),
    .io_in_addr(soundRomCache_1_io_in_addr),
    .io_in_dout(soundRomCache_1_io_in_dout),
    .io_in_wait_n(soundRomCache_1_io_in_wait_n),
    .io_in_valid(soundRomCache_1_io_in_valid),
    .io_out_rd(soundRomCache_1_io_out_rd),
    .io_out_addr(soundRomCache_1_io_out_addr),
    .io_out_dout(soundRomCache_1_io_out_dout),
    .io_out_wait_n(soundRomCache_1_io_out_wait_n),
    .io_out_valid(soundRomCache_1_io_out_valid)
  );
  ReadCache_3 layerRomCache_0 ( // @[MemSys.scala 149:19]
    .clock(layerRomCache_0_clock),
    .reset(layerRomCache_0_reset),
    .io_enable(layerRomCache_0_io_enable),
    .io_in_rd(layerRomCache_0_io_in_rd),
    .io_in_addr(layerRomCache_0_io_in_addr),
    .io_in_dout(layerRomCache_0_io_in_dout),
    .io_in_wait_n(layerRomCache_0_io_in_wait_n),
    .io_in_valid(layerRomCache_0_io_in_valid),
    .io_out_rd(layerRomCache_0_io_out_rd),
    .io_out_addr(layerRomCache_0_io_out_addr),
    .io_out_dout(layerRomCache_0_io_out_dout),
    .io_out_wait_n(layerRomCache_0_io_out_wait_n),
    .io_out_valid(layerRomCache_0_io_out_valid)
  );
  ReadCache_3 layerRomCache_1 ( // @[MemSys.scala 149:19]
    .clock(layerRomCache_1_clock),
    .reset(layerRomCache_1_reset),
    .io_enable(layerRomCache_1_io_enable),
    .io_in_rd(layerRomCache_1_io_in_rd),
    .io_in_addr(layerRomCache_1_io_in_addr),
    .io_in_dout(layerRomCache_1_io_in_dout),
    .io_in_wait_n(layerRomCache_1_io_in_wait_n),
    .io_in_valid(layerRomCache_1_io_in_valid),
    .io_out_rd(layerRomCache_1_io_out_rd),
    .io_out_addr(layerRomCache_1_io_out_addr),
    .io_out_dout(layerRomCache_1_io_out_dout),
    .io_out_wait_n(layerRomCache_1_io_out_wait_n),
    .io_out_valid(layerRomCache_1_io_out_valid)
  );
  ReadCache_3 layerRomCache_2 ( // @[MemSys.scala 149:19]
    .clock(layerRomCache_2_clock),
    .reset(layerRomCache_2_reset),
    .io_enable(layerRomCache_2_io_enable),
    .io_in_rd(layerRomCache_2_io_in_rd),
    .io_in_addr(layerRomCache_2_io_in_addr),
    .io_in_dout(layerRomCache_2_io_in_dout),
    .io_in_wait_n(layerRomCache_2_io_in_wait_n),
    .io_in_valid(layerRomCache_2_io_in_valid),
    .io_out_rd(layerRomCache_2_io_out_rd),
    .io_out_addr(layerRomCache_2_io_out_addr),
    .io_out_dout(layerRomCache_2_io_out_dout),
    .io_out_wait_n(layerRomCache_2_io_out_wait_n),
    .io_out_valid(layerRomCache_2_io_out_valid)
  );
  BurstMemArbiter ddrArbiter ( // @[MemSys.scala 164:26]
    .clock(ddrArbiter_clock),
    .reset(ddrArbiter_reset),
    .io_in_0_wr(ddrArbiter_io_in_0_wr),
    .io_in_0_addr(ddrArbiter_io_in_0_addr),
    .io_in_0_din(ddrArbiter_io_in_0_din),
    .io_in_0_burstDone(ddrArbiter_io_in_0_burstDone),
    .io_in_1_rd(ddrArbiter_io_in_1_rd),
    .io_in_1_addr(ddrArbiter_io_in_1_addr),
    .io_in_1_dout(ddrArbiter_io_in_1_dout),
    .io_in_1_wait_n(ddrArbiter_io_in_1_wait_n),
    .io_in_1_valid(ddrArbiter_io_in_1_valid),
    .io_in_1_burstDone(ddrArbiter_io_in_1_burstDone),
    .io_in_2_wr(ddrArbiter_io_in_2_wr),
    .io_in_2_addr(ddrArbiter_io_in_2_addr),
    .io_in_2_mask(ddrArbiter_io_in_2_mask),
    .io_in_2_din(ddrArbiter_io_in_2_din),
    .io_in_2_wait_n(ddrArbiter_io_in_2_wait_n),
    .io_in_3_rd(ddrArbiter_io_in_3_rd),
    .io_in_3_wr(ddrArbiter_io_in_3_wr),
    .io_in_3_addr(ddrArbiter_io_in_3_addr),
    .io_in_3_mask(ddrArbiter_io_in_3_mask),
    .io_in_3_din(ddrArbiter_io_in_3_din),
    .io_in_3_dout(ddrArbiter_io_in_3_dout),
    .io_in_3_wait_n(ddrArbiter_io_in_3_wait_n),
    .io_in_3_valid(ddrArbiter_io_in_3_valid),
    .io_in_3_burstLength(ddrArbiter_io_in_3_burstLength),
    .io_in_3_burstDone(ddrArbiter_io_in_3_burstDone),
    .io_in_4_rd(ddrArbiter_io_in_4_rd),
    .io_in_4_addr(ddrArbiter_io_in_4_addr),
    .io_in_4_dout(ddrArbiter_io_in_4_dout),
    .io_in_4_wait_n(ddrArbiter_io_in_4_wait_n),
    .io_in_4_valid(ddrArbiter_io_in_4_valid),
    .io_in_4_burstLength(ddrArbiter_io_in_4_burstLength),
    .io_in_4_burstDone(ddrArbiter_io_in_4_burstDone),
    .io_out_rd(ddrArbiter_io_out_rd),
    .io_out_wr(ddrArbiter_io_out_wr),
    .io_out_addr(ddrArbiter_io_out_addr),
    .io_out_mask(ddrArbiter_io_out_mask),
    .io_out_din(ddrArbiter_io_out_din),
    .io_out_dout(ddrArbiter_io_out_dout),
    .io_out_wait_n(ddrArbiter_io_out_wait_n),
    .io_out_valid(ddrArbiter_io_out_valid),
    .io_out_burstLength(ddrArbiter_io_out_burstLength),
    .io_out_burstDone(ddrArbiter_io_out_burstDone)
  );
  BurstMemArbiter_1 sdramArbiter ( // @[MemSys.scala 174:28]
    .clock(sdramArbiter_clock),
    .reset(sdramArbiter_reset),
    .io_in_0_wr(sdramArbiter_io_in_0_wr),
    .io_in_0_addr(sdramArbiter_io_in_0_addr),
    .io_in_0_din(sdramArbiter_io_in_0_din),
    .io_in_0_wait_n(sdramArbiter_io_in_0_wait_n),
    .io_in_0_burstDone(sdramArbiter_io_in_0_burstDone),
    .io_in_1_rd(sdramArbiter_io_in_1_rd),
    .io_in_1_addr(sdramArbiter_io_in_1_addr),
    .io_in_1_dout(sdramArbiter_io_in_1_dout),
    .io_in_1_wait_n(sdramArbiter_io_in_1_wait_n),
    .io_in_1_valid(sdramArbiter_io_in_1_valid),
    .io_in_2_rd(sdramArbiter_io_in_2_rd),
    .io_in_2_wr(sdramArbiter_io_in_2_wr),
    .io_in_2_addr(sdramArbiter_io_in_2_addr),
    .io_in_2_din(sdramArbiter_io_in_2_din),
    .io_in_2_dout(sdramArbiter_io_in_2_dout),
    .io_in_2_wait_n(sdramArbiter_io_in_2_wait_n),
    .io_in_2_valid(sdramArbiter_io_in_2_valid),
    .io_in_3_rd(sdramArbiter_io_in_3_rd),
    .io_in_3_addr(sdramArbiter_io_in_3_addr),
    .io_in_3_dout(sdramArbiter_io_in_3_dout),
    .io_in_3_wait_n(sdramArbiter_io_in_3_wait_n),
    .io_in_3_valid(sdramArbiter_io_in_3_valid),
    .io_in_4_rd(sdramArbiter_io_in_4_rd),
    .io_in_4_addr(sdramArbiter_io_in_4_addr),
    .io_in_4_dout(sdramArbiter_io_in_4_dout),
    .io_in_4_wait_n(sdramArbiter_io_in_4_wait_n),
    .io_in_4_valid(sdramArbiter_io_in_4_valid),
    .io_in_5_rd(sdramArbiter_io_in_5_rd),
    .io_in_5_addr(sdramArbiter_io_in_5_addr),
    .io_in_5_dout(sdramArbiter_io_in_5_dout),
    .io_in_5_wait_n(sdramArbiter_io_in_5_wait_n),
    .io_in_5_valid(sdramArbiter_io_in_5_valid),
    .io_in_6_rd(sdramArbiter_io_in_6_rd),
    .io_in_6_addr(sdramArbiter_io_in_6_addr),
    .io_in_6_dout(sdramArbiter_io_in_6_dout),
    .io_in_6_wait_n(sdramArbiter_io_in_6_wait_n),
    .io_in_6_valid(sdramArbiter_io_in_6_valid),
    .io_in_7_rd(sdramArbiter_io_in_7_rd),
    .io_in_7_addr(sdramArbiter_io_in_7_addr),
    .io_in_7_dout(sdramArbiter_io_in_7_dout),
    .io_in_7_wait_n(sdramArbiter_io_in_7_wait_n),
    .io_in_7_valid(sdramArbiter_io_in_7_valid),
    .io_out_rd(sdramArbiter_io_out_rd),
    .io_out_wr(sdramArbiter_io_out_wr),
    .io_out_addr(sdramArbiter_io_out_addr),
    .io_out_din(sdramArbiter_io_out_din),
    .io_out_dout(sdramArbiter_io_out_dout),
    .io_out_wait_n(sdramArbiter_io_out_wait_n),
    .io_out_valid(sdramArbiter_io_out_valid),
    .io_out_burstDone(sdramArbiter_io_out_burstDone)
  );
  AsyncMemArbiter nvramArbiter ( // @[MemSys.scala 187:28]
    .clock(nvramArbiter_clock),
    .reset(nvramArbiter_reset),
    .io_in_0_rd(nvramArbiter_io_in_0_rd),
    .io_in_0_wr(nvramArbiter_io_in_0_wr),
    .io_in_0_addr(nvramArbiter_io_in_0_addr),
    .io_in_0_din(nvramArbiter_io_in_0_din),
    .io_in_0_dout(nvramArbiter_io_in_0_dout),
    .io_in_0_wait_n(nvramArbiter_io_in_0_wait_n),
    .io_in_0_valid(nvramArbiter_io_in_0_valid),
    .io_in_1_rd(nvramArbiter_io_in_1_rd),
    .io_in_1_wr(nvramArbiter_io_in_1_wr),
    .io_in_1_addr(nvramArbiter_io_in_1_addr),
    .io_in_1_din(nvramArbiter_io_in_1_din),
    .io_in_1_dout(nvramArbiter_io_in_1_dout),
    .io_in_1_wait_n(nvramArbiter_io_in_1_wait_n),
    .io_in_1_valid(nvramArbiter_io_in_1_valid),
    .io_out_rd(nvramArbiter_io_out_rd),
    .io_out_wr(nvramArbiter_io_out_wr),
    .io_out_addr(nvramArbiter_io_out_addr),
    .io_out_din(nvramArbiter_io_out_din),
    .io_out_dout(nvramArbiter_io_out_dout),
    .io_out_wait_n(nvramArbiter_io_out_wait_n),
    .io_out_valid(nvramArbiter_io_out_valid)
  );
  assign io_prog_rom_wait_n = sdramDownloadBuffer_io_in_wait_n; // @[MemSys.scala 99:29]
  assign io_prog_nvram_dout = nvramArbiter_io_in_0_dout; // @[AsyncMemArbiter.scala 68:67]
  assign io_prog_nvram_wait_n = nvramArbiter_io_in_0_wait_n; // @[AsyncMemArbiter.scala 68:67]
  assign io_prog_nvram_valid = nvramArbiter_io_in_0_valid; // @[AsyncMemArbiter.scala 68:67]
  assign io_progRom_dout = progRomCache_io_in_dout; // @[MemSys.scala 117:22]
  assign io_progRom_wait_n = progRomCache_io_in_wait_n; // @[MemSys.scala 117:22]
  assign io_progRom_valid = progRomCache_io_in_valid; // @[MemSys.scala 117:22]
  assign io_eeprom_dout = nvramArbiter_io_in_1_dout; // @[AsyncMemArbiter.scala 68:67]
  assign io_eeprom_wait_n = nvramArbiter_io_in_1_wait_n; // @[AsyncMemArbiter.scala 68:67]
  assign io_eeprom_valid = nvramArbiter_io_in_1_valid; // @[AsyncMemArbiter.scala 68:67]
  assign io_soundRom_0_dout = soundRomCache_0_io_in_dout; // @[MemSys.scala 143:13]
  assign io_soundRom_0_wait_n = soundRomCache_0_io_in_wait_n; // @[MemSys.scala 143:13]
  assign io_soundRom_0_valid = soundRomCache_0_io_in_valid; // @[MemSys.scala 143:13]
  assign io_soundRom_1_dout = soundRomCache_1_io_in_dout; // @[MemSys.scala 143:13]
  assign io_soundRom_1_wait_n = soundRomCache_1_io_in_wait_n; // @[MemSys.scala 143:13]
  assign io_soundRom_1_valid = soundRomCache_1_io_in_valid; // @[MemSys.scala 143:13]
  assign io_layerTileRom_0_dout = layerRomCache_0_io_in_dout; // @[MemSys.scala 159:13]
  assign io_layerTileRom_0_wait_n = layerRomCache_0_io_in_wait_n; // @[MemSys.scala 159:13]
  assign io_layerTileRom_0_valid = layerRomCache_0_io_in_valid; // @[MemSys.scala 159:13]
  assign io_layerTileRom_1_dout = layerRomCache_1_io_in_dout; // @[MemSys.scala 159:13]
  assign io_layerTileRom_1_wait_n = layerRomCache_1_io_in_wait_n; // @[MemSys.scala 159:13]
  assign io_layerTileRom_1_valid = layerRomCache_1_io_in_valid; // @[MemSys.scala 159:13]
  assign io_layerTileRom_2_dout = layerRomCache_2_io_in_dout; // @[MemSys.scala 159:13]
  assign io_layerTileRom_2_wait_n = layerRomCache_2_io_in_wait_n; // @[MemSys.scala 159:13]
  assign io_layerTileRom_2_valid = layerRomCache_2_io_in_valid; // @[MemSys.scala 159:13]
  assign io_spriteTileRom_dout = ddrArbiter_io_in_4_dout; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign io_spriteTileRom_wait_n = ddrArbiter_io_in_4_wait_n; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign io_spriteTileRom_valid = ddrArbiter_io_in_4_valid; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign io_spriteTileRom_burstDone = ddrArbiter_io_in_4_burstDone; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign io_ddr_rd = ddrArbiter_io_out_rd; // @[MemSys.scala 171:5]
  assign io_ddr_wr = ddrArbiter_io_out_wr; // @[MemSys.scala 171:5]
  assign io_ddr_addr = ddrArbiter_io_out_addr; // @[MemSys.scala 171:5]
  assign io_ddr_mask = ddrArbiter_io_out_mask; // @[MemSys.scala 171:5]
  assign io_ddr_din = ddrArbiter_io_out_din; // @[MemSys.scala 171:5]
  assign io_ddr_burstLength = ddrArbiter_io_out_burstLength; // @[MemSys.scala 171:5]
  assign io_sdram_rd = sdramArbiter_io_out_rd; // @[MemSys.scala 184:5]
  assign io_sdram_wr = sdramArbiter_io_out_wr; // @[MemSys.scala 184:5]
  assign io_sdram_addr = sdramArbiter_io_out_addr; // @[MemSys.scala 184:5]
  assign io_sdram_din = sdramArbiter_io_out_din; // @[MemSys.scala 184:5]
  assign io_spriteFrameBuffer_dout = ddrArbiter_io_in_3_dout; // @[BurstMemArbiter.scala 68:67]
  assign io_spriteFrameBuffer_wait_n = ddrArbiter_io_in_3_wait_n; // @[BurstMemArbiter.scala 68:67]
  assign io_spriteFrameBuffer_valid = ddrArbiter_io_in_3_valid; // @[BurstMemArbiter.scala 68:67]
  assign io_spriteFrameBuffer_burstDone = ddrArbiter_io_in_3_burstDone; // @[BurstMemArbiter.scala 68:67]
  assign io_systemFrameBuffer_wait_n = ddrArbiter_io_in_2_wait_n; // @[BurstMemArbiter.scala 68:67]
  assign io_ready = io_ready_enableReg; // @[MemSys.scala 191:12]
  assign ddrDownloadBuffer_clock = clock;
  assign ddrDownloadBuffer_reset = reset;
  assign ddrDownloadBuffer_io_in_wr = io_prog_rom_wr; // @[MemSys.scala 88:27]
  assign ddrDownloadBuffer_io_in_addr = io_prog_rom_addr; // @[MemSys.scala 88:27]
  assign ddrDownloadBuffer_io_in_din = io_prog_rom_din; // @[MemSys.scala 88:27]
  assign ddrDownloadBuffer_io_out_burstDone = ddrArbiter_io_in_0_burstDone; // @[BurstMemIO.scala 156:19 BurstMemArbiter.scala 68:67]
  assign sdramDownloadBuffer_clock = clock;
  assign sdramDownloadBuffer_reset = reset;
  assign sdramDownloadBuffer_io_in_wr = copyDma_io_out_wr; // @[MemSys.scala 104:18]
  assign sdramDownloadBuffer_io_in_addr = copyDma_io_out_addr; // @[MemSys.scala 104:18]
  assign sdramDownloadBuffer_io_in_din = copyDma_io_out_din; // @[MemSys.scala 104:18]
  assign sdramDownloadBuffer_io_out_wait_n = sdramArbiter_io_in_0_wait_n; // @[BurstMemIO.scala 156:19 BurstMemArbiter.scala 68:67]
  assign sdramDownloadBuffer_io_out_burstDone = sdramArbiter_io_in_0_burstDone; // @[BurstMemIO.scala 156:19 BurstMemArbiter.scala 68:67]
  assign copyDma_clock = clock;
  assign copyDma_reset = reset;
  assign copyDma_io_start = ~io_ready & io_prog_done; // @[MemSys.scala 103:33]
  assign copyDma_io_in_dout = ddrArbiter_io_in_1_dout; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign copyDma_io_in_wait_n = ddrArbiter_io_in_1_wait_n; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign copyDma_io_in_valid = ddrArbiter_io_in_1_valid; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign copyDma_io_in_burstDone = ddrArbiter_io_in_1_burstDone; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign copyDma_io_out_wait_n = sdramDownloadBuffer_io_in_wait_n; // @[MemSys.scala 104:18]
  assign progRomCache_clock = clock;
  assign progRomCache_reset = reset;
  assign progRomCache_io_enable = io_ready; // @[MemSys.scala 116:26]
  assign progRomCache_io_in_rd = io_progRom_rd; // @[MemSys.scala 117:22]
  assign progRomCache_io_in_addr = io_progRom_addr; // @[MemSys.scala 117:22]
  assign progRomCache_io_out_dout = sdramArbiter_io_in_1_dout; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign progRomCache_io_out_wait_n = sdramArbiter_io_in_1_wait_n; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign progRomCache_io_out_valid = sdramArbiter_io_in_1_valid; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign eepromCache_clock = clock;
  assign eepromCache_reset = reset;
  assign eepromCache_io_enable = io_ready; // @[MemSys.scala 129:25]
  assign eepromCache_io_in_rd = nvramArbiter_io_out_rd; // @[MemSys.scala 188:50]
  assign eepromCache_io_in_wr = nvramArbiter_io_out_wr; // @[MemSys.scala 188:50]
  assign eepromCache_io_in_addr = nvramArbiter_io_out_addr; // @[MemSys.scala 188:50]
  assign eepromCache_io_in_din = nvramArbiter_io_out_din; // @[MemSys.scala 188:50]
  assign eepromCache_io_out_dout = sdramArbiter_io_in_2_dout; // @[BurstMemIO.scala 269:19 BurstMemArbiter.scala 68:67]
  assign eepromCache_io_out_wait_n = sdramArbiter_io_in_2_wait_n; // @[BurstMemIO.scala 269:19 BurstMemArbiter.scala 68:67]
  assign eepromCache_io_out_valid = sdramArbiter_io_in_2_valid; // @[BurstMemIO.scala 269:19 BurstMemArbiter.scala 68:67]
  assign soundRomCache_0_clock = clock;
  assign soundRomCache_0_reset = reset;
  assign soundRomCache_0_io_enable = io_ready; // @[MemSys.scala 142:17]
  assign soundRomCache_0_io_in_rd = io_soundRom_0_rd; // @[MemSys.scala 143:13]
  assign soundRomCache_0_io_in_addr = io_soundRom_0_addr; // @[MemSys.scala 143:13]
  assign soundRomCache_0_io_out_dout = sdramArbiter_io_in_3_dout; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign soundRomCache_0_io_out_wait_n = sdramArbiter_io_in_3_wait_n; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign soundRomCache_0_io_out_valid = sdramArbiter_io_in_3_valid; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign soundRomCache_1_clock = clock;
  assign soundRomCache_1_reset = reset;
  assign soundRomCache_1_io_enable = io_ready; // @[MemSys.scala 142:17]
  assign soundRomCache_1_io_in_rd = io_soundRom_1_rd; // @[MemSys.scala 143:13]
  assign soundRomCache_1_io_in_addr = io_soundRom_1_addr; // @[MemSys.scala 143:13]
  assign soundRomCache_1_io_out_dout = sdramArbiter_io_in_4_dout; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign soundRomCache_1_io_out_wait_n = sdramArbiter_io_in_4_wait_n; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign soundRomCache_1_io_out_valid = sdramArbiter_io_in_4_valid; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign layerRomCache_0_clock = clock;
  assign layerRomCache_0_reset = reset;
  assign layerRomCache_0_io_enable = io_ready; // @[MemSys.scala 158:17]
  assign layerRomCache_0_io_in_rd = io_layerTileRom_0_rd; // @[MemSys.scala 159:13]
  assign layerRomCache_0_io_in_addr = io_layerTileRom_0_addr; // @[MemSys.scala 159:13]
  assign layerRomCache_0_io_out_dout = sdramArbiter_io_in_5_dout; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign layerRomCache_0_io_out_wait_n = sdramArbiter_io_in_5_wait_n; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign layerRomCache_0_io_out_valid = sdramArbiter_io_in_5_valid; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign layerRomCache_1_clock = clock;
  assign layerRomCache_1_reset = reset;
  assign layerRomCache_1_io_enable = io_ready; // @[MemSys.scala 158:17]
  assign layerRomCache_1_io_in_rd = io_layerTileRom_1_rd; // @[MemSys.scala 159:13]
  assign layerRomCache_1_io_in_addr = io_layerTileRom_1_addr; // @[MemSys.scala 159:13]
  assign layerRomCache_1_io_out_dout = sdramArbiter_io_in_6_dout; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign layerRomCache_1_io_out_wait_n = sdramArbiter_io_in_6_wait_n; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign layerRomCache_1_io_out_valid = sdramArbiter_io_in_6_valid; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign layerRomCache_2_clock = clock;
  assign layerRomCache_2_reset = reset;
  assign layerRomCache_2_io_enable = io_ready; // @[MemSys.scala 158:17]
  assign layerRomCache_2_io_in_rd = io_layerTileRom_2_rd; // @[MemSys.scala 159:13]
  assign layerRomCache_2_io_in_addr = io_layerTileRom_2_addr; // @[MemSys.scala 159:13]
  assign layerRomCache_2_io_out_dout = sdramArbiter_io_in_7_dout; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign layerRomCache_2_io_out_wait_n = sdramArbiter_io_in_7_wait_n; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign layerRomCache_2_io_out_valid = sdramArbiter_io_in_7_valid; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign ddrArbiter_clock = clock;
  assign ddrArbiter_reset = reset;
  assign ddrArbiter_io_in_0_wr = ddrDownloadBuffer_io_out_wr; // @[BurstMemIO.scala 180:19 181:12]
  assign ddrArbiter_io_in_0_addr = ddrDownloadBuffer_io_out_addr + 32'h30000000; // @[MemSys.scala 166:40]
  assign ddrArbiter_io_in_0_din = ddrDownloadBuffer_io_out_din; // @[BurstMemIO.scala 180:19 187:13]
  assign ddrArbiter_io_in_1_rd = copyDma_io_in_rd; // @[BurstMemIO.scala 89:19 90:12]
  assign ddrArbiter_io_in_1_addr = copyDma_io_in_addr + 32'h30000000; // @[MemSys.scala 167:29]
  assign ddrArbiter_io_in_2_wr = io_systemFrameBuffer_wr; // @[BurstMemArbiter.scala 68:67]
  assign ddrArbiter_io_in_2_addr = io_systemFrameBuffer_addr; // @[BurstMemArbiter.scala 68:67]
  assign ddrArbiter_io_in_2_mask = io_systemFrameBuffer_mask; // @[BurstMemArbiter.scala 68:67]
  assign ddrArbiter_io_in_2_din = io_systemFrameBuffer_din; // @[BurstMemArbiter.scala 68:67]
  assign ddrArbiter_io_in_3_rd = io_spriteFrameBuffer_rd; // @[BurstMemArbiter.scala 68:67]
  assign ddrArbiter_io_in_3_wr = io_spriteFrameBuffer_wr; // @[BurstMemArbiter.scala 68:67]
  assign ddrArbiter_io_in_3_addr = io_spriteFrameBuffer_addr; // @[BurstMemArbiter.scala 68:67]
  assign ddrArbiter_io_in_3_mask = io_spriteFrameBuffer_mask; // @[BurstMemArbiter.scala 68:67]
  assign ddrArbiter_io_in_3_din = io_spriteFrameBuffer_din; // @[BurstMemArbiter.scala 68:67]
  assign ddrArbiter_io_in_3_burstLength = io_spriteFrameBuffer_burstLength; // @[BurstMemArbiter.scala 68:67]
  assign ddrArbiter_io_in_4_rd = io_spriteTileRom_rd; // @[BurstMemIO.scala 89:19 90:12]
  assign ddrArbiter_io_in_4_addr = _mem_T_5 + 32'h30000000; // @[MemSys.scala 170:65]
  assign ddrArbiter_io_in_4_burstLength = io_spriteTileRom_burstLength; // @[BurstMemIO.scala 89:19 91:21]
  assign ddrArbiter_io_out_dout = io_ddr_dout; // @[MemSys.scala 171:5]
  assign ddrArbiter_io_out_wait_n = io_ddr_wait_n; // @[MemSys.scala 171:5]
  assign ddrArbiter_io_out_valid = io_ddr_valid; // @[MemSys.scala 171:5]
  assign ddrArbiter_io_out_burstDone = io_ddr_burstDone; // @[MemSys.scala 171:5]
  assign sdramArbiter_clock = clock;
  assign sdramArbiter_reset = reset;
  assign sdramArbiter_io_in_0_wr = sdramDownloadBuffer_io_out_wr; // @[BurstMemIO.scala 156:19 158:12]
  assign sdramArbiter_io_in_0_addr = sdramDownloadBuffer_io_out_addr; // @[BurstMemIO.scala 156:19 162:14]
  assign sdramArbiter_io_in_0_din = sdramDownloadBuffer_io_out_din; // @[BurstMemIO.scala 156:19 164:13]
  assign sdramArbiter_io_in_1_rd = progRomCache_io_out_rd; // @[BurstMemIO.scala 89:19 90:12]
  assign sdramArbiter_io_in_1_addr = _mem_T_8[24:0]; // @[BurstMemArbiter.scala 68:67]
  assign sdramArbiter_io_in_2_rd = eepromCache_io_out_rd; // @[BurstMemIO.scala 269:19 270:12]
  assign sdramArbiter_io_in_2_wr = eepromCache_io_out_wr; // @[BurstMemIO.scala 269:19 271:12]
  assign sdramArbiter_io_in_2_addr = _mem_T_11[24:0]; // @[BurstMemArbiter.scala 68:67]
  assign sdramArbiter_io_in_2_din = eepromCache_io_out_din; // @[BurstMemIO.scala 269:19 278:13]
  assign sdramArbiter_io_in_3_rd = soundRomCache_0_io_out_rd; // @[BurstMemIO.scala 89:19 90:12]
  assign sdramArbiter_io_in_3_addr = _mem_T_13[24:0]; // @[BurstMemArbiter.scala 68:67]
  assign sdramArbiter_io_in_4_rd = soundRomCache_1_io_out_rd; // @[BurstMemIO.scala 89:19 90:12]
  assign sdramArbiter_io_in_4_addr = _mem_T_15[24:0]; // @[BurstMemArbiter.scala 68:67]
  assign sdramArbiter_io_in_5_rd = layerRomCache_0_io_out_rd; // @[BurstMemIO.scala 89:19 90:12]
  assign sdramArbiter_io_in_5_addr = _mem_T_17[24:0]; // @[BurstMemArbiter.scala 68:67]
  assign sdramArbiter_io_in_6_rd = layerRomCache_1_io_out_rd; // @[BurstMemIO.scala 89:19 90:12]
  assign sdramArbiter_io_in_6_addr = _mem_T_19[24:0]; // @[BurstMemArbiter.scala 68:67]
  assign sdramArbiter_io_in_7_rd = layerRomCache_2_io_out_rd; // @[BurstMemIO.scala 89:19 90:12]
  assign sdramArbiter_io_in_7_addr = _mem_T_21[24:0]; // @[BurstMemArbiter.scala 68:67]
  assign sdramArbiter_io_out_dout = io_sdram_dout; // @[MemSys.scala 184:5]
  assign sdramArbiter_io_out_wait_n = io_sdram_wait_n; // @[MemSys.scala 184:5]
  assign sdramArbiter_io_out_valid = io_sdram_valid; // @[MemSys.scala 184:5]
  assign sdramArbiter_io_out_burstDone = io_sdram_burstDone; // @[MemSys.scala 184:5]
  assign nvramArbiter_clock = clock;
  assign nvramArbiter_reset = reset;
  assign nvramArbiter_io_in_0_rd = io_prog_nvram_rd; // @[AsyncMemArbiter.scala 68:67]
  assign nvramArbiter_io_in_0_wr = io_prog_nvram_wr; // @[AsyncMemArbiter.scala 68:67]
  assign nvramArbiter_io_in_0_addr = io_prog_nvram_addr[6:0]; // @[AsyncMemArbiter.scala 68:67]
  assign nvramArbiter_io_in_0_din = io_prog_nvram_din; // @[AsyncMemArbiter.scala 68:67]
  assign nvramArbiter_io_in_1_rd = io_eeprom_rd; // @[AsyncMemArbiter.scala 68:67]
  assign nvramArbiter_io_in_1_wr = io_eeprom_wr; // @[AsyncMemArbiter.scala 68:67]
  assign nvramArbiter_io_in_1_addr = io_eeprom_addr; // @[AsyncMemArbiter.scala 68:67]
  assign nvramArbiter_io_in_1_din = io_eeprom_din; // @[AsyncMemArbiter.scala 68:67]
  assign nvramArbiter_io_out_dout = eepromCache_io_in_dout; // @[MemSys.scala 188:50]
  assign nvramArbiter_io_out_wait_n = eepromCache_io_in_wait_n; // @[MemSys.scala 188:50]
  assign nvramArbiter_io_out_valid = eepromCache_io_in_valid; // @[MemSys.scala 188:50]
  always @(posedge clock) begin
    io_ready_REG <= copyDma_io_busy; // @[Util.scala 165:45]
    if (reset) begin // @[Util.scala 218:28]
      io_ready_enableReg <= 1'h0; // @[Util.scala 218:28]
    end else begin
      io_ready_enableReg <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_ready_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_ready_enableReg = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegisterFile_1(
  input         clock,
  input         io_mem_wr,
  input  [2:0]  io_mem_addr,
  input  [15:0] io_mem_din,
  output [15:0] io_regs_0,
  output [15:0] io_regs_1,
  output [15:0] io_regs_2,
  output [15:0] io_regs_3,
  output [15:0] io_regs_4,
  output [15:0] io_regs_5
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] regs_0; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_1; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_2; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_3; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_4; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_5; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_6; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_7; // @[RegisterFile.scala 56:17]
  wire [15:0] _GEN_1 = 3'h1 == io_mem_addr ? regs_1 : regs_0; // @[]
  wire [15:0] _GEN_2 = 3'h2 == io_mem_addr ? regs_2 : _GEN_1; // @[]
  wire [15:0] _GEN_3 = 3'h3 == io_mem_addr ? regs_3 : _GEN_2; // @[]
  wire [15:0] _GEN_4 = 3'h4 == io_mem_addr ? regs_4 : _GEN_3; // @[]
  wire [15:0] _GEN_5 = 3'h5 == io_mem_addr ? regs_5 : _GEN_4; // @[]
  wire [15:0] _GEN_6 = 3'h6 == io_mem_addr ? regs_6 : _GEN_5; // @[]
  wire [15:0] _GEN_7 = 3'h7 == io_mem_addr ? regs_7 : _GEN_6; // @[]
  wire [7:0] bytes_0 = io_mem_wr ? io_mem_din[7:0] : _GEN_7[7:0]; // @[RegisterFile.scala 62:28 66:{39,50}]
  wire [7:0] bytes_1 = io_mem_wr ? io_mem_din[15:8] : _GEN_7[15:8]; // @[RegisterFile.scala 62:28 66:{39,50}]
  wire [15:0] _regs_T = {bytes_1,bytes_0}; // @[RegisterFile.scala 70:17]
  assign io_regs_0 = regs_0; // @[RegisterFile.scala 74:11]
  assign io_regs_1 = regs_1; // @[RegisterFile.scala 74:11]
  assign io_regs_2 = regs_2; // @[RegisterFile.scala 74:11]
  assign io_regs_3 = regs_3; // @[RegisterFile.scala 74:11]
  assign io_regs_4 = regs_4; // @[RegisterFile.scala 74:11]
  assign io_regs_5 = regs_5; // @[RegisterFile.scala 74:11]
  always @(posedge clock) begin
    if (3'h0 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_0 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h1 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_1 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h2 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_2 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h3 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_3 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h4 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_4 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h5 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_5 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h6 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_6 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h7 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_7 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module VideoTiming(
  input        clock,
  input        reset,
  input  [8:0] io_display_x,
  input  [8:0] io_display_y,
  input  [8:0] io_frontPorch_x,
  input  [8:0] io_frontPorch_y,
  input  [8:0] io_retrace_x,
  input  [8:0] io_retrace_y,
  input  [3:0] io_offset_x,
  input  [3:0] io_offset_y,
  output       io_timing_clockEnable,
  output       io_timing_displayEnable,
  output [8:0] io_timing_pos_x,
  output [8:0] io_timing_pos_y,
  output       io_timing_hSync,
  output       io_timing_vSync,
  output       io_timing_hBlank,
  output       io_timing_vBlank
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] clockDivWrap_value; // @[Counter.scala 40:34]
  wire  clockDivWrap_wrap_wrap = clockDivWrap_value == 2'h3; // @[Counter.scala 45:24]
  wire [1:0] _clockDivWrap_wrap_value_T_1 = clockDivWrap_value + 2'h1; // @[Counter.scala 46:22]
  reg [8:0] x; // @[Counter.scala 40:34]
  wire  wrap_wrap = x == 9'h1bf; // @[Counter.scala 45:24]
  wire [8:0] _wrap_value_T_1 = x + 9'h1; // @[Counter.scala 46:22]
  wire  xWrap = clockDivWrap_wrap_wrap & wrap_wrap; // @[Counter.scala 86:{48,55}]
  wire  _T = clockDivWrap_wrap_wrap & xWrap; // @[VideoTiming.scala 89:72]
  reg [8:0] y; // @[Counter.scala 40:34]
  wire  wrap_wrap_1 = y == 9'h10f; // @[Counter.scala 45:24]
  wire [8:0] _wrap_value_T_3 = y + 9'h1; // @[Counter.scala 46:22]
  wire [9:0] _GEN_14 = {{6{io_offset_x[3]}},io_offset_x}; // @[VideoTiming.scala 92:39]
  wire [9:0] _hBeginDisplay_T_3 = 10'sh1c0 + $signed(_GEN_14); // @[VideoTiming.scala 92:54]
  wire [9:0] _GEN_15 = {{1'd0}, io_display_x}; // @[VideoTiming.scala 92:61]
  wire [9:0] _hBeginDisplay_T_5 = _hBeginDisplay_T_3 - _GEN_15; // @[VideoTiming.scala 92:61]
  wire [9:0] _GEN_16 = {{1'd0}, io_frontPorch_x}; // @[VideoTiming.scala 92:76]
  wire [9:0] _hBeginDisplay_T_7 = _hBeginDisplay_T_5 - _GEN_16; // @[VideoTiming.scala 92:76]
  wire [9:0] _GEN_17 = {{1'd0}, io_retrace_x}; // @[VideoTiming.scala 92:94]
  wire [9:0] hBeginDisplay = _hBeginDisplay_T_7 - _GEN_17; // @[VideoTiming.scala 92:94]
  wire [9:0] _hEndDisplay_T_5 = _hBeginDisplay_T_3 - _GEN_16; // @[VideoTiming.scala 93:59]
  wire [9:0] hEndDisplay = _hEndDisplay_T_5 - _GEN_17; // @[VideoTiming.scala 93:77]
  wire [8:0] hBeginSync = 9'h1c0 - io_retrace_x; // @[VideoTiming.scala 94:35]
  wire [9:0] _GEN_21 = {{6{io_offset_y[3]}},io_offset_y}; // @[VideoTiming.scala 98:40]
  wire [9:0] _vBeginDisplay_T_3 = 10'sh110 + $signed(_GEN_21); // @[VideoTiming.scala 98:55]
  wire [9:0] _GEN_22 = {{1'd0}, io_display_y}; // @[VideoTiming.scala 98:62]
  wire [9:0] _vBeginDisplay_T_5 = _vBeginDisplay_T_3 - _GEN_22; // @[VideoTiming.scala 98:62]
  wire [9:0] _GEN_23 = {{1'd0}, io_frontPorch_y}; // @[VideoTiming.scala 98:77]
  wire [9:0] _vBeginDisplay_T_7 = _vBeginDisplay_T_5 - _GEN_23; // @[VideoTiming.scala 98:77]
  wire [9:0] _GEN_24 = {{1'd0}, io_retrace_y}; // @[VideoTiming.scala 98:95]
  wire [9:0] vBeginDisplay = _vBeginDisplay_T_7 - _GEN_24; // @[VideoTiming.scala 98:95]
  wire [9:0] _vEndDisplay_T_5 = _vBeginDisplay_T_3 - _GEN_23; // @[VideoTiming.scala 99:60]
  wire [9:0] vEndDisplay = _vEndDisplay_T_5 - _GEN_24; // @[VideoTiming.scala 99:78]
  wire [8:0] vBeginSync = 9'h110 - io_retrace_y; // @[VideoTiming.scala 100:36]
  wire [9:0] _GEN_28 = {{1'd0}, x}; // @[VideoTiming.scala 104:21]
  wire [9:0] pos_x = _GEN_28 - hBeginDisplay; // @[VideoTiming.scala 104:21]
  wire [9:0] _GEN_29 = {{1'd0}, y}; // @[VideoTiming.scala 104:40]
  wire [9:0] pos_y = _GEN_29 - vBeginDisplay; // @[VideoTiming.scala 104:40]
  wire  hBlank = _GEN_28 < hBeginDisplay | _GEN_28 >= hEndDisplay; // @[VideoTiming.scala 111:34]
  wire  vBlank = _GEN_29 < vBeginDisplay | _GEN_29 >= vEndDisplay; // @[VideoTiming.scala 112:34]
  assign io_timing_clockEnable = clockDivWrap_value == 2'h3; // @[Counter.scala 45:24]
  assign io_timing_displayEnable = ~(hBlank | vBlank); // @[VideoTiming.scala 116:30]
  assign io_timing_pos_x = pos_x[8:0]; // @[VideoTiming.scala 117:17]
  assign io_timing_pos_y = pos_y[8:0]; // @[VideoTiming.scala 117:17]
  assign io_timing_hSync = x >= hBeginSync & x < 9'h1c0; // @[VideoTiming.scala 107:31]
  assign io_timing_vSync = y >= vBeginSync & y < 9'h110; // @[VideoTiming.scala 108:31]
  assign io_timing_hBlank = _GEN_28 < hBeginDisplay | _GEN_28 >= hEndDisplay; // @[VideoTiming.scala 111:34]
  assign io_timing_vBlank = _GEN_29 < vBeginDisplay | _GEN_29 >= vEndDisplay; // @[VideoTiming.scala 112:34]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 40:34]
      clockDivWrap_value <= 2'h0; // @[Counter.scala 40:34]
    end else begin
      clockDivWrap_value <= _clockDivWrap_wrap_value_T_1;
    end
    if (reset) begin // @[Counter.scala 40:34]
      x <= 9'h0; // @[Counter.scala 40:34]
    end else if (clockDivWrap_wrap_wrap) begin // @[Counter.scala 86:48]
      if (wrap_wrap) begin // @[Counter.scala 48:20]
        x <= 9'h0; // @[Counter.scala 48:28]
      end else begin
        x <= _wrap_value_T_1; // @[Counter.scala 46:13]
      end
    end
    if (reset) begin // @[Counter.scala 40:34]
      y <= 9'h0; // @[Counter.scala 40:34]
    end else if (_T) begin // @[Counter.scala 86:48]
      if (wrap_wrap_1) begin // @[Counter.scala 48:20]
        y <= 9'h0; // @[Counter.scala 48:28]
      end else begin
        y <= _wrap_value_T_3; // @[Counter.scala 46:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  clockDivWrap_value = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  x = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  y = _RAND_2[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module VideoTiming_1(
  input        clock,
  input        reset,
  input  [8:0] io_display_x,
  input  [8:0] io_display_y,
  input  [8:0] io_frontPorch_x,
  input  [8:0] io_frontPorch_y,
  input  [8:0] io_retrace_x,
  input  [8:0] io_retrace_y,
  input  [3:0] io_offset_x,
  input  [3:0] io_offset_y,
  output       io_timing_clockEnable,
  output       io_timing_displayEnable,
  output [8:0] io_timing_pos_x,
  output [8:0] io_timing_pos_y,
  output       io_timing_hSync,
  output       io_timing_vSync,
  output       io_timing_hBlank,
  output       io_timing_vBlank
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] clockDivWrap_value; // @[Counter.scala 40:34]
  wire  clockDivWrap_wrap_wrap = clockDivWrap_value == 2'h3; // @[Counter.scala 45:24]
  wire [1:0] _clockDivWrap_wrap_value_T_1 = clockDivWrap_value + 2'h1; // @[Counter.scala 46:22]
  reg [8:0] x; // @[Counter.scala 40:34]
  wire  wrap_wrap = x == 9'h1bc; // @[Counter.scala 45:24]
  wire [8:0] _wrap_value_T_1 = x + 9'h1; // @[Counter.scala 46:22]
  wire  xWrap = clockDivWrap_wrap_wrap & wrap_wrap; // @[Counter.scala 86:{48,55}]
  wire  _T = clockDivWrap_wrap_wrap & xWrap; // @[VideoTiming.scala 89:72]
  reg [8:0] y; // @[Counter.scala 40:34]
  wire  wrap_wrap_1 = y == 9'h105; // @[Counter.scala 45:24]
  wire [8:0] _wrap_value_T_3 = y + 9'h1; // @[Counter.scala 46:22]
  wire [9:0] _GEN_14 = {{6{io_offset_x[3]}},io_offset_x}; // @[VideoTiming.scala 92:39]
  wire [9:0] _hBeginDisplay_T_3 = 10'sh1bd + $signed(_GEN_14); // @[VideoTiming.scala 92:54]
  wire [9:0] _GEN_15 = {{1'd0}, io_display_x}; // @[VideoTiming.scala 92:61]
  wire [9:0] _hBeginDisplay_T_5 = _hBeginDisplay_T_3 - _GEN_15; // @[VideoTiming.scala 92:61]
  wire [9:0] _GEN_16 = {{1'd0}, io_frontPorch_x}; // @[VideoTiming.scala 92:76]
  wire [9:0] _hBeginDisplay_T_7 = _hBeginDisplay_T_5 - _GEN_16; // @[VideoTiming.scala 92:76]
  wire [9:0] _GEN_17 = {{1'd0}, io_retrace_x}; // @[VideoTiming.scala 92:94]
  wire [9:0] hBeginDisplay = _hBeginDisplay_T_7 - _GEN_17; // @[VideoTiming.scala 92:94]
  wire [9:0] _hEndDisplay_T_5 = _hBeginDisplay_T_3 - _GEN_16; // @[VideoTiming.scala 93:59]
  wire [9:0] hEndDisplay = _hEndDisplay_T_5 - _GEN_17; // @[VideoTiming.scala 93:77]
  wire [8:0] hBeginSync = 9'h1bd - io_retrace_x; // @[VideoTiming.scala 94:35]
  wire [9:0] _GEN_21 = {{6{io_offset_y[3]}},io_offset_y}; // @[VideoTiming.scala 98:40]
  wire [9:0] _vBeginDisplay_T_3 = 10'sh106 + $signed(_GEN_21); // @[VideoTiming.scala 98:55]
  wire [9:0] _GEN_22 = {{1'd0}, io_display_y}; // @[VideoTiming.scala 98:62]
  wire [9:0] _vBeginDisplay_T_5 = _vBeginDisplay_T_3 - _GEN_22; // @[VideoTiming.scala 98:62]
  wire [9:0] _GEN_23 = {{1'd0}, io_frontPorch_y}; // @[VideoTiming.scala 98:77]
  wire [9:0] _vBeginDisplay_T_7 = _vBeginDisplay_T_5 - _GEN_23; // @[VideoTiming.scala 98:77]
  wire [9:0] _GEN_24 = {{1'd0}, io_retrace_y}; // @[VideoTiming.scala 98:95]
  wire [9:0] vBeginDisplay = _vBeginDisplay_T_7 - _GEN_24; // @[VideoTiming.scala 98:95]
  wire [9:0] _vEndDisplay_T_5 = _vBeginDisplay_T_3 - _GEN_23; // @[VideoTiming.scala 99:60]
  wire [9:0] vEndDisplay = _vEndDisplay_T_5 - _GEN_24; // @[VideoTiming.scala 99:78]
  wire [8:0] vBeginSync = 9'h106 - io_retrace_y; // @[VideoTiming.scala 100:36]
  wire [9:0] _GEN_28 = {{1'd0}, x}; // @[VideoTiming.scala 104:21]
  wire [9:0] pos_x = _GEN_28 - hBeginDisplay; // @[VideoTiming.scala 104:21]
  wire [9:0] _GEN_29 = {{1'd0}, y}; // @[VideoTiming.scala 104:40]
  wire [9:0] pos_y = _GEN_29 - vBeginDisplay; // @[VideoTiming.scala 104:40]
  wire  hBlank = _GEN_28 < hBeginDisplay | _GEN_28 >= hEndDisplay; // @[VideoTiming.scala 111:34]
  wire  vBlank = _GEN_29 < vBeginDisplay | _GEN_29 >= vEndDisplay; // @[VideoTiming.scala 112:34]
  assign io_timing_clockEnable = clockDivWrap_value == 2'h3; // @[Counter.scala 45:24]
  assign io_timing_displayEnable = ~(hBlank | vBlank); // @[VideoTiming.scala 116:30]
  assign io_timing_pos_x = pos_x[8:0]; // @[VideoTiming.scala 117:17]
  assign io_timing_pos_y = pos_y[8:0]; // @[VideoTiming.scala 117:17]
  assign io_timing_hSync = x >= hBeginSync & x < 9'h1bd; // @[VideoTiming.scala 107:31]
  assign io_timing_vSync = y >= vBeginSync & y < 9'h106; // @[VideoTiming.scala 108:31]
  assign io_timing_hBlank = _GEN_28 < hBeginDisplay | _GEN_28 >= hEndDisplay; // @[VideoTiming.scala 111:34]
  assign io_timing_vBlank = _GEN_29 < vBeginDisplay | _GEN_29 >= vEndDisplay; // @[VideoTiming.scala 112:34]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 40:34]
      clockDivWrap_value <= 2'h0; // @[Counter.scala 40:34]
    end else begin
      clockDivWrap_value <= _clockDivWrap_wrap_value_T_1;
    end
    if (reset) begin // @[Counter.scala 40:34]
      x <= 9'h0; // @[Counter.scala 40:34]
    end else if (clockDivWrap_wrap_wrap) begin // @[Counter.scala 86:48]
      if (wrap_wrap) begin // @[Counter.scala 48:20]
        x <= 9'h0; // @[Counter.scala 48:28]
      end else begin
        x <= _wrap_value_T_1; // @[Counter.scala 46:13]
      end
    end
    if (reset) begin // @[Counter.scala 40:34]
      y <= 9'h0; // @[Counter.scala 40:34]
    end else if (_T) begin // @[Counter.scala 86:48]
      if (wrap_wrap_1) begin // @[Counter.scala 48:20]
        y <= 9'h0; // @[Counter.scala 48:28]
      end else begin
        y <= _wrap_value_T_3; // @[Counter.scala 46:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  clockDivWrap_value = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  x = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  y = _RAND_2[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module VideoSys(
  input         clock,
  input         reset,
  input         io_videoClock,
  input         io_videoReset,
  input         io_prog_video_wr,
  input  [26:0] io_prog_video_addr,
  input  [15:0] io_prog_video_din,
  input         io_prog_done,
  input  [3:0]  io_options_offset_x,
  input  [3:0]  io_options_offset_y,
  input         io_options_compatibility,
  output        io_video_clockEnable,
  output        io_video_displayEnable,
  output [8:0]  io_video_pos_x,
  output [8:0]  io_video_pos_y,
  output        io_video_hSync,
  output        io_video_vSync,
  output        io_video_hBlank,
  output        io_video_vBlank,
  output [8:0]  io_video_regs_size_x,
  output [8:0]  io_video_regs_size_y,
  output [8:0]  io_video_regs_frontPorch_x,
  output [8:0]  io_video_regs_frontPorch_y,
  output [8:0]  io_video_regs_retrace_x,
  output [8:0]  io_video_regs_retrace_y,
  output        io_video_changeMode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire  videoRegs_clock; // @[VideoSys.scala 66:25]
  wire  videoRegs_io_mem_wr; // @[VideoSys.scala 66:25]
  wire [2:0] videoRegs_io_mem_addr; // @[VideoSys.scala 66:25]
  wire [15:0] videoRegs_io_mem_din; // @[VideoSys.scala 66:25]
  wire [15:0] videoRegs_io_regs_0; // @[VideoSys.scala 66:25]
  wire [15:0] videoRegs_io_regs_1; // @[VideoSys.scala 66:25]
  wire [15:0] videoRegs_io_regs_2; // @[VideoSys.scala 66:25]
  wire [15:0] videoRegs_io_regs_3; // @[VideoSys.scala 66:25]
  wire [15:0] videoRegs_io_regs_4; // @[VideoSys.scala 66:25]
  wire [15:0] videoRegs_io_regs_5; // @[VideoSys.scala 66:25]
  wire  timing_originalVideoTiming_clock; // @[VideoSys.scala 74:37]
  wire  timing_originalVideoTiming_reset; // @[VideoSys.scala 74:37]
  wire [8:0] timing_originalVideoTiming_io_display_x; // @[VideoSys.scala 74:37]
  wire [8:0] timing_originalVideoTiming_io_display_y; // @[VideoSys.scala 74:37]
  wire [8:0] timing_originalVideoTiming_io_frontPorch_x; // @[VideoSys.scala 74:37]
  wire [8:0] timing_originalVideoTiming_io_frontPorch_y; // @[VideoSys.scala 74:37]
  wire [8:0] timing_originalVideoTiming_io_retrace_x; // @[VideoSys.scala 74:37]
  wire [8:0] timing_originalVideoTiming_io_retrace_y; // @[VideoSys.scala 74:37]
  wire [3:0] timing_originalVideoTiming_io_offset_x; // @[VideoSys.scala 74:37]
  wire [3:0] timing_originalVideoTiming_io_offset_y; // @[VideoSys.scala 74:37]
  wire  timing_originalVideoTiming_io_timing_clockEnable; // @[VideoSys.scala 74:37]
  wire  timing_originalVideoTiming_io_timing_displayEnable; // @[VideoSys.scala 74:37]
  wire [8:0] timing_originalVideoTiming_io_timing_pos_x; // @[VideoSys.scala 74:37]
  wire [8:0] timing_originalVideoTiming_io_timing_pos_y; // @[VideoSys.scala 74:37]
  wire  timing_originalVideoTiming_io_timing_hSync; // @[VideoSys.scala 74:37]
  wire  timing_originalVideoTiming_io_timing_vSync; // @[VideoSys.scala 74:37]
  wire  timing_originalVideoTiming_io_timing_hBlank; // @[VideoSys.scala 74:37]
  wire  timing_originalVideoTiming_io_timing_vBlank; // @[VideoSys.scala 74:37]
  wire  timing_compatibilityVideoTiming_clock; // @[VideoSys.scala 80:42]
  wire  timing_compatibilityVideoTiming_reset; // @[VideoSys.scala 80:42]
  wire [8:0] timing_compatibilityVideoTiming_io_display_x; // @[VideoSys.scala 80:42]
  wire [8:0] timing_compatibilityVideoTiming_io_display_y; // @[VideoSys.scala 80:42]
  wire [8:0] timing_compatibilityVideoTiming_io_frontPorch_x; // @[VideoSys.scala 80:42]
  wire [8:0] timing_compatibilityVideoTiming_io_frontPorch_y; // @[VideoSys.scala 80:42]
  wire [8:0] timing_compatibilityVideoTiming_io_retrace_x; // @[VideoSys.scala 80:42]
  wire [8:0] timing_compatibilityVideoTiming_io_retrace_y; // @[VideoSys.scala 80:42]
  wire [3:0] timing_compatibilityVideoTiming_io_offset_x; // @[VideoSys.scala 80:42]
  wire [3:0] timing_compatibilityVideoTiming_io_offset_y; // @[VideoSys.scala 80:42]
  wire  timing_compatibilityVideoTiming_io_timing_clockEnable; // @[VideoSys.scala 80:42]
  wire  timing_compatibilityVideoTiming_io_timing_displayEnable; // @[VideoSys.scala 80:42]
  wire [8:0] timing_compatibilityVideoTiming_io_timing_pos_x; // @[VideoSys.scala 80:42]
  wire [8:0] timing_compatibilityVideoTiming_io_timing_pos_y; // @[VideoSys.scala 80:42]
  wire  timing_compatibilityVideoTiming_io_timing_hSync; // @[VideoSys.scala 80:42]
  wire  timing_compatibilityVideoTiming_io_timing_vSync; // @[VideoSys.scala 80:42]
  wire  timing_compatibilityVideoTiming_io_timing_hBlank; // @[VideoSys.scala 80:42]
  wire  timing_compatibilityVideoTiming_io_timing_vBlank; // @[VideoSys.scala 80:42]
  reg [3:0] timing_originalVideoTiming_io_offset_r_x; // @[Reg.scala 19:16]
  reg [3:0] timing_originalVideoTiming_io_offset_r_y; // @[Reg.scala 19:16]
  reg [3:0] timing_compatibilityVideoTiming_io_offset_r_x; // @[Reg.scala 19:16]
  reg [3:0] timing_compatibilityVideoTiming_io_offset_r_y; // @[Reg.scala 19:16]
  wire  _timing_latchReg_T = timing_originalVideoTiming_io_timing_vBlank &
    timing_compatibilityVideoTiming_io_timing_vBlank; // @[VideoSys.scala 93:93]
  reg  timing_latchReg; // @[Reg.scala 19:16]
  reg  timing_clockEnable; // @[VideoSys.scala 99:12]
  reg  timing_displayEnable; // @[VideoSys.scala 99:12]
  reg [8:0] timing_pos_x; // @[VideoSys.scala 99:12]
  reg [8:0] timing_pos_y; // @[VideoSys.scala 99:12]
  reg  timing_hSync; // @[VideoSys.scala 99:12]
  reg  timing_vSync; // @[VideoSys.scala 99:12]
  reg  timing_hBlank; // @[VideoSys.scala 99:12]
  reg  timing_vBlank; // @[VideoSys.scala 99:12]
  wire [8:0] io_video_regs_regs_size_vec_x = videoRegs_io_regs_0[8:0]; // @[VideoRegs.scala 92:31]
  wire [8:0] io_video_regs_regs_size_vec_y = videoRegs_io_regs_1[8:0]; // @[VideoRegs.scala 92:46]
  wire [8:0] io_video_regs_regs_frontPorch_vec_x = videoRegs_io_regs_2[8:0]; // @[VideoRegs.scala 93:37]
  wire [8:0] io_video_regs_regs_frontPorch_vec_y = videoRegs_io_regs_3[8:0]; // @[VideoRegs.scala 93:52]
  wire [8:0] io_video_regs_regs_retrace_vec_x = videoRegs_io_regs_4[8:0] + 9'h8; // @[VideoRegs.scala 94:41]
  wire [8:0] io_video_regs_regs_retrace_vec_y = videoRegs_io_regs_5[8:0] + 9'h1; // @[VideoRegs.scala 94:62]
  reg [8:0] io_video_regs_r_size_x; // @[Reg.scala 35:20]
  reg [8:0] io_video_regs_r_size_y; // @[Reg.scala 35:20]
  reg [8:0] io_video_regs_r_frontPorch_x; // @[Reg.scala 35:20]
  reg [8:0] io_video_regs_r_frontPorch_y; // @[Reg.scala 35:20]
  reg [8:0] io_video_regs_r_retrace_x; // @[Reg.scala 35:20]
  reg [8:0] io_video_regs_r_retrace_y; // @[Reg.scala 35:20]
  reg  io_video_changeMode_REG; // @[VideoSys.scala 111:77]
  RegisterFile_1 videoRegs ( // @[VideoSys.scala 66:25]
    .clock(videoRegs_clock),
    .io_mem_wr(videoRegs_io_mem_wr),
    .io_mem_addr(videoRegs_io_mem_addr),
    .io_mem_din(videoRegs_io_mem_din),
    .io_regs_0(videoRegs_io_regs_0),
    .io_regs_1(videoRegs_io_regs_1),
    .io_regs_2(videoRegs_io_regs_2),
    .io_regs_3(videoRegs_io_regs_3),
    .io_regs_4(videoRegs_io_regs_4),
    .io_regs_5(videoRegs_io_regs_5)
  );
  VideoTiming timing_originalVideoTiming ( // @[VideoSys.scala 74:37]
    .clock(timing_originalVideoTiming_clock),
    .reset(timing_originalVideoTiming_reset),
    .io_display_x(timing_originalVideoTiming_io_display_x),
    .io_display_y(timing_originalVideoTiming_io_display_y),
    .io_frontPorch_x(timing_originalVideoTiming_io_frontPorch_x),
    .io_frontPorch_y(timing_originalVideoTiming_io_frontPorch_y),
    .io_retrace_x(timing_originalVideoTiming_io_retrace_x),
    .io_retrace_y(timing_originalVideoTiming_io_retrace_y),
    .io_offset_x(timing_originalVideoTiming_io_offset_x),
    .io_offset_y(timing_originalVideoTiming_io_offset_y),
    .io_timing_clockEnable(timing_originalVideoTiming_io_timing_clockEnable),
    .io_timing_displayEnable(timing_originalVideoTiming_io_timing_displayEnable),
    .io_timing_pos_x(timing_originalVideoTiming_io_timing_pos_x),
    .io_timing_pos_y(timing_originalVideoTiming_io_timing_pos_y),
    .io_timing_hSync(timing_originalVideoTiming_io_timing_hSync),
    .io_timing_vSync(timing_originalVideoTiming_io_timing_vSync),
    .io_timing_hBlank(timing_originalVideoTiming_io_timing_hBlank),
    .io_timing_vBlank(timing_originalVideoTiming_io_timing_vBlank)
  );
  VideoTiming_1 timing_compatibilityVideoTiming ( // @[VideoSys.scala 80:42]
    .clock(timing_compatibilityVideoTiming_clock),
    .reset(timing_compatibilityVideoTiming_reset),
    .io_display_x(timing_compatibilityVideoTiming_io_display_x),
    .io_display_y(timing_compatibilityVideoTiming_io_display_y),
    .io_frontPorch_x(timing_compatibilityVideoTiming_io_frontPorch_x),
    .io_frontPorch_y(timing_compatibilityVideoTiming_io_frontPorch_y),
    .io_retrace_x(timing_compatibilityVideoTiming_io_retrace_x),
    .io_retrace_y(timing_compatibilityVideoTiming_io_retrace_y),
    .io_offset_x(timing_compatibilityVideoTiming_io_offset_x),
    .io_offset_y(timing_compatibilityVideoTiming_io_offset_y),
    .io_timing_clockEnable(timing_compatibilityVideoTiming_io_timing_clockEnable),
    .io_timing_displayEnable(timing_compatibilityVideoTiming_io_timing_displayEnable),
    .io_timing_pos_x(timing_compatibilityVideoTiming_io_timing_pos_x),
    .io_timing_pos_y(timing_compatibilityVideoTiming_io_timing_pos_y),
    .io_timing_hSync(timing_compatibilityVideoTiming_io_timing_hSync),
    .io_timing_vSync(timing_compatibilityVideoTiming_io_timing_vSync),
    .io_timing_hBlank(timing_compatibilityVideoTiming_io_timing_hBlank),
    .io_timing_vBlank(timing_compatibilityVideoTiming_io_timing_vBlank)
  );
  assign io_video_clockEnable = timing_clockEnable; // @[VideoSys.scala 103:24]
  assign io_video_displayEnable = timing_displayEnable; // @[VideoSys.scala 104:26]
  assign io_video_pos_x = timing_pos_x; // @[VideoSys.scala 105:16]
  assign io_video_pos_y = timing_pos_y; // @[VideoSys.scala 105:16]
  assign io_video_hSync = timing_hSync; // @[VideoSys.scala 106:18]
  assign io_video_vSync = timing_vSync; // @[VideoSys.scala 107:18]
  assign io_video_hBlank = timing_hBlank; // @[VideoSys.scala 108:19]
  assign io_video_vBlank = timing_vBlank; // @[VideoSys.scala 109:19]
  assign io_video_regs_size_x = io_video_regs_r_size_x; // @[VideoSys.scala 110:17]
  assign io_video_regs_size_y = io_video_regs_r_size_y; // @[VideoSys.scala 110:17]
  assign io_video_regs_frontPorch_x = io_video_regs_r_frontPorch_x; // @[VideoSys.scala 110:17]
  assign io_video_regs_frontPorch_y = io_video_regs_r_frontPorch_y; // @[VideoSys.scala 110:17]
  assign io_video_regs_retrace_x = io_video_regs_r_retrace_x; // @[VideoSys.scala 110:17]
  assign io_video_regs_retrace_y = io_video_regs_r_retrace_y; // @[VideoSys.scala 110:17]
  assign io_video_changeMode = io_prog_done | io_options_compatibility ^ io_video_changeMode_REG; // @[VideoSys.scala 111:39]
  assign videoRegs_clock = clock;
  assign videoRegs_io_mem_wr = io_prog_video_wr; // @[AsyncMemIO.scala 236:19 237:12]
  assign videoRegs_io_mem_addr = io_prog_video_addr[3:1]; // @[VideoSys.scala 67:20]
  assign videoRegs_io_mem_din = {io_prog_video_din[7:0],io_prog_video_din[15:8]}; // @[Util.scala 114:49]
  assign timing_originalVideoTiming_clock = io_videoClock;
  assign timing_originalVideoTiming_reset = io_videoReset;
  assign timing_originalVideoTiming_io_display_x = io_video_regs_size_x; // @[VideoSys.scala 75:36]
  assign timing_originalVideoTiming_io_display_y = io_video_regs_size_y; // @[VideoSys.scala 75:36]
  assign timing_originalVideoTiming_io_frontPorch_x = io_video_regs_frontPorch_x; // @[VideoSys.scala 76:39]
  assign timing_originalVideoTiming_io_frontPorch_y = io_video_regs_frontPorch_y; // @[VideoSys.scala 76:39]
  assign timing_originalVideoTiming_io_retrace_x = io_video_regs_retrace_x; // @[VideoSys.scala 77:36]
  assign timing_originalVideoTiming_io_retrace_y = io_video_regs_retrace_y; // @[VideoSys.scala 77:36]
  assign timing_originalVideoTiming_io_offset_x = timing_originalVideoTiming_io_offset_r_x; // @[VideoSys.scala 88:35]
  assign timing_originalVideoTiming_io_offset_y = timing_originalVideoTiming_io_offset_r_y; // @[VideoSys.scala 88:35]
  assign timing_compatibilityVideoTiming_clock = io_videoClock;
  assign timing_compatibilityVideoTiming_reset = io_videoReset;
  assign timing_compatibilityVideoTiming_io_display_x = io_video_regs_size_x; // @[VideoSys.scala 81:41]
  assign timing_compatibilityVideoTiming_io_display_y = io_video_regs_size_y; // @[VideoSys.scala 81:41]
  assign timing_compatibilityVideoTiming_io_frontPorch_x = io_video_regs_frontPorch_x; // @[VideoSys.scala 82:44]
  assign timing_compatibilityVideoTiming_io_frontPorch_y = io_video_regs_frontPorch_y; // @[VideoSys.scala 82:44]
  assign timing_compatibilityVideoTiming_io_retrace_x = io_video_regs_retrace_x; // @[VideoSys.scala 83:41]
  assign timing_compatibilityVideoTiming_io_retrace_y = io_video_regs_retrace_y; // @[VideoSys.scala 83:41]
  assign timing_compatibilityVideoTiming_io_offset_x = timing_compatibilityVideoTiming_io_offset_r_x; // @[VideoSys.scala 89:40]
  assign timing_compatibilityVideoTiming_io_offset_y = timing_compatibilityVideoTiming_io_offset_r_y; // @[VideoSys.scala 89:40]
  always @(posedge io_videoClock) begin
    if (timing_originalVideoTiming_io_timing_vSync) begin // @[Reg.scala 20:18]
      timing_originalVideoTiming_io_offset_r_x <= io_options_offset_x; // @[Reg.scala 20:22]
    end
    if (timing_originalVideoTiming_io_timing_vSync) begin // @[Reg.scala 20:18]
      timing_originalVideoTiming_io_offset_r_y <= io_options_offset_y; // @[Reg.scala 20:22]
    end
    if (timing_compatibilityVideoTiming_io_timing_vSync) begin // @[Reg.scala 20:18]
      timing_compatibilityVideoTiming_io_offset_r_x <= io_options_offset_x; // @[Reg.scala 20:22]
    end
    if (timing_compatibilityVideoTiming_io_timing_vSync) begin // @[Reg.scala 20:18]
      timing_compatibilityVideoTiming_io_offset_r_y <= io_options_offset_y; // @[Reg.scala 20:22]
    end
    if (_timing_latchReg_T) begin // @[Reg.scala 20:18]
      timing_latchReg <= io_options_compatibility; // @[Reg.scala 20:22]
    end
    if (timing_latchReg) begin // @[VideoSys.scala 96:21]
      timing_clockEnable <= timing_compatibilityVideoTiming_io_timing_clockEnable;
    end else begin
      timing_clockEnable <= timing_originalVideoTiming_io_timing_clockEnable;
    end
    if (timing_latchReg) begin // @[VideoSys.scala 96:21]
      timing_displayEnable <= timing_compatibilityVideoTiming_io_timing_displayEnable;
    end else begin
      timing_displayEnable <= timing_originalVideoTiming_io_timing_displayEnable;
    end
    if (timing_latchReg) begin // @[VideoSys.scala 96:21]
      timing_pos_x <= timing_compatibilityVideoTiming_io_timing_pos_x;
    end else begin
      timing_pos_x <= timing_originalVideoTiming_io_timing_pos_x;
    end
    if (timing_latchReg) begin // @[VideoSys.scala 96:21]
      timing_pos_y <= timing_compatibilityVideoTiming_io_timing_pos_y;
    end else begin
      timing_pos_y <= timing_originalVideoTiming_io_timing_pos_y;
    end
    if (timing_latchReg) begin // @[VideoSys.scala 96:21]
      timing_hSync <= timing_compatibilityVideoTiming_io_timing_hSync;
    end else begin
      timing_hSync <= timing_originalVideoTiming_io_timing_hSync;
    end
    if (timing_latchReg) begin // @[VideoSys.scala 96:21]
      timing_vSync <= timing_compatibilityVideoTiming_io_timing_vSync;
    end else begin
      timing_vSync <= timing_originalVideoTiming_io_timing_vSync;
    end
    if (timing_latchReg) begin // @[VideoSys.scala 96:21]
      timing_hBlank <= timing_compatibilityVideoTiming_io_timing_hBlank;
    end else begin
      timing_hBlank <= timing_originalVideoTiming_io_timing_hBlank;
    end
    if (timing_latchReg) begin // @[VideoSys.scala 96:21]
      timing_vBlank <= timing_compatibilityVideoTiming_io_timing_vBlank;
    end else begin
      timing_vBlank <= timing_originalVideoTiming_io_timing_vBlank;
    end
  end
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      io_video_regs_r_size_x <= 9'h140; // @[Reg.scala 35:20]
    end else if (io_prog_done) begin // @[Reg.scala 36:18]
      io_video_regs_r_size_x <= io_video_regs_regs_size_vec_x; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      io_video_regs_r_size_y <= 9'hf0; // @[Reg.scala 35:20]
    end else if (io_prog_done) begin // @[Reg.scala 36:18]
      io_video_regs_r_size_y <= io_video_regs_regs_size_vec_y; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      io_video_regs_r_frontPorch_x <= 9'h24; // @[Reg.scala 35:20]
    end else if (io_prog_done) begin // @[Reg.scala 36:18]
      io_video_regs_r_frontPorch_x <= io_video_regs_regs_frontPorch_vec_x; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      io_video_regs_r_frontPorch_y <= 9'hc; // @[Reg.scala 35:20]
    end else if (io_prog_done) begin // @[Reg.scala 36:18]
      io_video_regs_r_frontPorch_y <= io_video_regs_regs_frontPorch_vec_y; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      io_video_regs_r_retrace_x <= 9'h1c; // @[Reg.scala 35:20]
    end else if (io_prog_done) begin // @[Reg.scala 36:18]
      io_video_regs_r_retrace_x <= io_video_regs_regs_retrace_vec_x; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      io_video_regs_r_retrace_y <= 9'h3; // @[Reg.scala 35:20]
    end else if (io_prog_done) begin // @[Reg.scala 36:18]
      io_video_regs_r_retrace_y <= io_video_regs_regs_retrace_vec_y; // @[Reg.scala 36:22]
    end
    io_video_changeMode_REG <= io_options_compatibility; // @[VideoSys.scala 111:77]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  timing_originalVideoTiming_io_offset_r_x = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  timing_originalVideoTiming_io_offset_r_y = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  timing_compatibilityVideoTiming_io_offset_r_x = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  timing_compatibilityVideoTiming_io_offset_r_y = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  timing_latchReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  timing_clockEnable = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  timing_displayEnable = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  timing_pos_x = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  timing_pos_y = _RAND_8[8:0];
  _RAND_9 = {1{`RANDOM}};
  timing_hSync = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  timing_vSync = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  timing_hBlank = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  timing_vBlank = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  io_video_regs_r_size_x = _RAND_13[8:0];
  _RAND_14 = {1{`RANDOM}};
  io_video_regs_r_size_y = _RAND_14[8:0];
  _RAND_15 = {1{`RANDOM}};
  io_video_regs_r_frontPorch_x = _RAND_15[8:0];
  _RAND_16 = {1{`RANDOM}};
  io_video_regs_r_frontPorch_y = _RAND_16[8:0];
  _RAND_17 = {1{`RANDOM}};
  io_video_regs_r_retrace_x = _RAND_17[8:0];
  _RAND_18 = {1{`RANDOM}};
  io_video_regs_r_retrace_y = _RAND_18[8:0];
  _RAND_19 = {1{`RANDOM}};
  io_video_changeMode_REG = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CPU(
  input         clock,
  input         reset,
  input         io_halt,
  output        io_as,
  output        io_rw,
  output        io_uds,
  output        io_lds,
  input         io_dtack,
  input         io_vpa,
  input  [2:0]  io_ipl,
  output [2:0]  io_fc,
  output [22:0] io_addr,
  input  [15:0] io_din,
  output [15:0] io_dout
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  cpu_clk; // @[CPU.scala 118:19]
  wire  cpu_enPhi1; // @[CPU.scala 118:19]
  wire  cpu_enPhi2; // @[CPU.scala 118:19]
  wire  cpu_extReset; // @[CPU.scala 118:19]
  wire  cpu_pwrUp; // @[CPU.scala 118:19]
  wire  cpu_HALTn; // @[CPU.scala 118:19]
  wire  cpu_ASn; // @[CPU.scala 118:19]
  wire  cpu_eRWn; // @[CPU.scala 118:19]
  wire  cpu_UDSn; // @[CPU.scala 118:19]
  wire  cpu_LDSn; // @[CPU.scala 118:19]
  wire  cpu_DTACKn; // @[CPU.scala 118:19]
  wire  cpu_BERRn; // @[CPU.scala 118:19]
  wire  cpu_E; // @[CPU.scala 118:19]
  wire  cpu_VPAn; // @[CPU.scala 118:19]
  wire  cpu_VMAn; // @[CPU.scala 118:19]
  wire  cpu_BRn; // @[CPU.scala 118:19]
  wire  cpu_BGn; // @[CPU.scala 118:19]
  wire  cpu_BGACKn; // @[CPU.scala 118:19]
  wire  cpu_IPL0n; // @[CPU.scala 118:19]
  wire  cpu_IPL1n; // @[CPU.scala 118:19]
  wire  cpu_IPL2n; // @[CPU.scala 118:19]
  wire  cpu_FC0; // @[CPU.scala 118:19]
  wire  cpu_FC1; // @[CPU.scala 118:19]
  wire  cpu_FC2; // @[CPU.scala 118:19]
  wire [22:0] cpu_eab; // @[CPU.scala 118:19]
  wire [15:0] cpu_iEdb; // @[CPU.scala 118:19]
  wire [15:0] cpu_oEdb; // @[CPU.scala 118:19]
  reg  phi1_value; // @[Counter.scala 40:34]
  wire  _phi1_wrap_value_T_1 = phi1_value + 1'h1; // @[Counter.scala 46:22]
  reg  phi2; // @[Reg.scala 19:16]
  wire [1:0] io_fc_hi = {cpu_FC2,cpu_FC1}; // @[Cat.scala 33:92]
  fx68k cpu ( // @[CPU.scala 118:19]
    .clk(cpu_clk),
    .enPhi1(cpu_enPhi1),
    .enPhi2(cpu_enPhi2),
    .extReset(cpu_extReset),
    .pwrUp(cpu_pwrUp),
    .HALTn(cpu_HALTn),
    .ASn(cpu_ASn),
    .eRWn(cpu_eRWn),
    .UDSn(cpu_UDSn),
    .LDSn(cpu_LDSn),
    .DTACKn(cpu_DTACKn),
    .BERRn(cpu_BERRn),
    .E(cpu_E),
    .VPAn(cpu_VPAn),
    .VMAn(cpu_VMAn),
    .BRn(cpu_BRn),
    .BGn(cpu_BGn),
    .BGACKn(cpu_BGACKn),
    .IPL0n(cpu_IPL0n),
    .IPL1n(cpu_IPL1n),
    .IPL2n(cpu_IPL2n),
    .FC0(cpu_FC0),
    .FC1(cpu_FC1),
    .FC2(cpu_FC2),
    .eab(cpu_eab),
    .iEdb(cpu_iEdb),
    .oEdb(cpu_oEdb)
  );
  assign io_as = ~cpu_ASn; // @[CPU.scala 125:12]
  assign io_rw = cpu_eRWn; // @[CPU.scala 126:9]
  assign io_uds = ~cpu_UDSn; // @[CPU.scala 127:13]
  assign io_lds = ~cpu_LDSn; // @[CPU.scala 128:13]
  assign io_fc = {io_fc_hi,cpu_FC0}; // @[Cat.scala 33:92]
  assign io_addr = cpu_eab; // @[CPU.scala 138:11]
  assign io_dout = cpu_oEdb; // @[CPU.scala 140:11]
  assign cpu_clk = clock; // @[CPU.scala 119:23]
  assign cpu_enPhi1 = phi1_value; // @[Counter.scala 86:17]
  assign cpu_enPhi2 = phi2; // @[CPU.scala 121:17]
  assign cpu_extReset = reset; // @[CPU.scala 122:28]
  assign cpu_pwrUp = reset; // @[CPU.scala 123:25]
  assign cpu_HALTn = ~io_halt; // @[CPU.scala 124:19]
  assign cpu_DTACKn = ~io_dtack; // @[CPU.scala 129:20]
  assign cpu_BERRn = 1'h1; // @[CPU.scala 130:16]
  assign cpu_VPAn = ~io_vpa; // @[CPU.scala 133:18]
  assign cpu_BRn = 1'h1; // @[CPU.scala 131:14]
  assign cpu_BGACKn = 1'h1; // @[CPU.scala 132:17]
  assign cpu_IPL0n = ~io_ipl[0]; // @[CPU.scala 134:19]
  assign cpu_IPL1n = ~io_ipl[1]; // @[CPU.scala 135:19]
  assign cpu_IPL2n = ~io_ipl[2]; // @[CPU.scala 136:19]
  assign cpu_iEdb = io_din; // @[CPU.scala 139:15]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 40:34]
      phi1_value <= 1'h0; // @[Counter.scala 40:34]
    end else begin
      phi1_value <= _phi1_wrap_value_T_1;
    end
    phi2 <= phi1_value; // @[Reg.scala 19:16 20:{18,22}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phi1_value = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  phi2 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EEPROM(
  input         clock,
  input         reset,
  output        io_mem_rd,
  output        io_mem_wr,
  output [6:0]  io_mem_addr,
  output [15:0] io_mem_din,
  input  [15:0] io_mem_dout,
  input         io_mem_wait_n,
  input         io_mem_valid,
  input         io_serial_cs,
  input         io_serial_sck,
  input         io_serial_sdi,
  output        io_serial_sdo
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] stateReg; // @[EEPROM.scala 65:25]
  reg [16:0] counterReg; // @[EEPROM.scala 68:27]
  reg [5:0] addrReg; // @[EEPROM.scala 69:20]
  reg [15:0] dataReg; // @[EEPROM.scala 70:20]
  reg [1:0] opcodeReg; // @[EEPROM.scala 71:22]
  reg  serialReg; // @[EEPROM.scala 72:26]
  reg  writeAllReg; // @[EEPROM.scala 73:28]
  reg  writeEnableReg; // @[EEPROM.scala 74:31]
  reg  sckRising_REG; // @[Util.scala 158:44]
  wire  sckRising = io_serial_sck & ~sckRising_REG; // @[Util.scala 158:33]
  wire  done = counterReg[0]; // @[EEPROM.scala 80:24]
  wire  read = opcodeReg == 2'h2; // @[EEPROM.scala 81:24]
  wire  write = opcodeReg == 2'h1 & writeEnableReg; // @[EEPROM.scala 82:33]
  wire  erase = opcodeReg == 2'h3 & writeEnableReg; // @[EEPROM.scala 83:33]
  wire  _writeAll_T = opcodeReg == 2'h0; // @[EEPROM.scala 84:28]
  wire  writeAll = opcodeReg == 2'h0 & addrReg[4:3] == 2'h1 & writeEnableReg; // @[EEPROM.scala 84:61]
  wire  eraseAll = _writeAll_T & addrReg[4:3] == 2'h2 & writeEnableReg; // @[EEPROM.scala 85:61]
  wire  enableWrite = _writeAll_T & addrReg[4:3] == 2'h3; // @[EEPROM.scala 86:39]
  wire  disableWrite = _writeAll_T & addrReg[4:3] == 2'h0; // @[EEPROM.scala 87:40]
  wire [16:0] _GEN_0 = (stateReg == 3'h2 | stateReg == 3'h6 | stateReg == 3'h7) & sckRising ? {{1'd0}, counterReg[16:1]}
     : counterReg; // @[EEPROM.scala 90:112 91:16 68:27]
  wire [2:0] _GEN_2 = sckRising & io_serial_sdi ? 3'h2 : stateReg; // @[EEPROM.scala 111:{40,51} 95:12]
  wire [8:0] data = {opcodeReg,addrReg,io_serial_sdi}; // @[EEPROM.scala 117:41]
  wire  _GEN_3 = disableWrite ? 1'h0 : writeEnableReg; // @[EEPROM.scala 147:36 148:28 74:31]
  wire  _GEN_5 = enableWrite | _GEN_3; // @[EEPROM.scala 144:35 145:28]
  wire [5:0] _GEN_7 = eraseAll ? 6'h0 : data[5:0]; // @[EEPROM.scala 123:17 140:32 141:21]
  wire  _GEN_8 = eraseAll | writeAllReg; // @[EEPROM.scala 140:32 142:25 73:28]
  wire [2:0] _GEN_9 = eraseAll ? 3'h5 : 3'h0; // @[EEPROM.scala 140:32 143:22]
  wire  _GEN_10 = eraseAll ? writeEnableReg : _GEN_5; // @[EEPROM.scala 140:32 74:31]
  wire [16:0] _GEN_11 = writeAll ? 17'h8000 : _GEN_0; // @[EEPROM.scala 135:32 136:24]
  wire [5:0] _GEN_12 = writeAll ? 6'h0 : _GEN_7; // @[EEPROM.scala 135:32 137:21]
  wire  _GEN_13 = writeAll | _GEN_8; // @[EEPROM.scala 135:32 138:25]
  wire [2:0] _GEN_14 = writeAll ? 3'h6 : _GEN_9; // @[EEPROM.scala 135:32 139:22]
  wire  _GEN_15 = writeAll ? writeEnableReg : _GEN_10; // @[EEPROM.scala 135:32 74:31]
  wire [2:0] _GEN_16 = erase ? 3'h5 : _GEN_14; // @[EEPROM.scala 133:29 134:22]
  wire [16:0] _GEN_17 = erase ? _GEN_0 : _GEN_11; // @[EEPROM.scala 133:29]
  wire [5:0] _GEN_18 = erase ? data[5:0] : _GEN_12; // @[EEPROM.scala 123:17 133:29]
  wire  _GEN_19 = erase ? writeAllReg : _GEN_13; // @[EEPROM.scala 133:29 73:28]
  wire  _GEN_20 = erase ? writeEnableReg : _GEN_15; // @[EEPROM.scala 133:29 74:31]
  wire [16:0] _GEN_21 = write ? 17'h8000 : _GEN_17; // @[EEPROM.scala 130:29 131:24]
  wire [2:0] _GEN_22 = write ? 3'h6 : _GEN_16; // @[EEPROM.scala 130:29 132:22]
  wire [5:0] _GEN_23 = write ? data[5:0] : _GEN_18; // @[EEPROM.scala 123:17 130:29]
  wire  _GEN_24 = write ? writeAllReg : _GEN_19; // @[EEPROM.scala 130:29 73:28]
  wire  _GEN_25 = write ? writeEnableReg : _GEN_20; // @[EEPROM.scala 130:29 74:31]
  wire [16:0] _GEN_26 = read ? 17'h10000 : _GEN_21; // @[EEPROM.scala 126:22 127:24]
  wire  _GEN_27 = read ? 1'h0 : serialReg; // @[EEPROM.scala 126:22 128:23 72:26]
  wire [2:0] _GEN_28 = read ? 3'h3 : _GEN_22; // @[EEPROM.scala 126:22 129:22]
  wire [5:0] _GEN_29 = read ? data[5:0] : _GEN_23; // @[EEPROM.scala 123:17 126:22]
  wire  _GEN_30 = read ? writeAllReg : _GEN_24; // @[EEPROM.scala 126:22 73:28]
  wire  _GEN_31 = read ? writeEnableReg : _GEN_25; // @[EEPROM.scala 126:22 74:31]
  wire [16:0] _GEN_32 = done ? _GEN_26 : _GEN_0; // @[EEPROM.scala 125:20]
  wire  _GEN_33 = done ? _GEN_27 : serialReg; // @[EEPROM.scala 125:20 72:26]
  wire [2:0] _GEN_34 = done ? _GEN_28 : stateReg; // @[EEPROM.scala 125:20 95:12]
  wire [5:0] _GEN_35 = done ? _GEN_29 : data[5:0]; // @[EEPROM.scala 123:17 125:20]
  wire  _GEN_36 = done ? _GEN_30 : writeAllReg; // @[EEPROM.scala 125:20 73:28]
  wire  _GEN_37 = done ? _GEN_31 : writeEnableReg; // @[EEPROM.scala 125:20 74:31]
  wire [16:0] _GEN_40 = sckRising ? _GEN_32 : _GEN_0; // @[EEPROM.scala 116:23]
  wire  _GEN_41 = sckRising ? _GEN_33 : serialReg; // @[EEPROM.scala 116:23 72:26]
  wire [2:0] _GEN_42 = sckRising ? _GEN_34 : stateReg; // @[EEPROM.scala 116:23 95:12]
  wire  _GEN_43 = sckRising ? _GEN_36 : writeAllReg; // @[EEPROM.scala 116:23 73:28]
  wire  _GEN_44 = sckRising ? _GEN_37 : writeEnableReg; // @[EEPROM.scala 116:23 74:31]
  wire [2:0] _GEN_45 = io_mem_wait_n ? 3'h4 : stateReg; // @[EEPROM.scala 162:33 163:18 95:12]
  wire [15:0] _GEN_46 = io_mem_valid ? io_mem_dout : dataReg; // @[EEPROM.scala 159:26 160:17 70:20]
  wire [2:0] _GEN_47 = io_mem_valid ? 3'h7 : _GEN_45; // @[EEPROM.scala 159:26 161:18]
  wire [2:0] _GEN_48 = io_mem_valid ? 3'h7 : stateReg; // @[EEPROM.scala 169:26 171:18 95:12]
  wire [5:0] _addrReg_T_2 = addrReg + 6'h1; // @[EEPROM.scala 178:28]
  wire [2:0] _GEN_49 = ~writeAllReg | &addrReg ? 3'h0 : stateReg; // @[EEPROM.scala 179:{44,55} 95:12]
  wire [5:0] _GEN_50 = io_mem_wait_n ? _addrReg_T_2 : addrReg; // @[EEPROM.scala 177:27 178:17 69:20]
  wire [2:0] _GEN_51 = io_mem_wait_n ? _GEN_49 : stateReg; // @[EEPROM.scala 177:27 95:12]
  wire [16:0] _dataReg_T = {dataReg,io_serial_sdi}; // @[EEPROM.scala 187:28]
  wire [2:0] _GEN_52 = done ? 3'h5 : stateReg; // @[EEPROM.scala 188:{20,31} 95:12]
  wire  _GEN_53 = sckRising ? 1'h0 : serialReg; // @[EEPROM.scala 185:23 186:19 72:26]
  wire [16:0] _GEN_54 = sckRising ? _dataReg_T : {{1'd0}, dataReg}; // @[EEPROM.scala 185:23 187:17 70:20]
  wire [2:0] _GEN_55 = sckRising ? _GEN_52 : stateReg; // @[EEPROM.scala 185:23 95:12]
  wire [16:0] _dataReg_T_1 = {dataReg,1'h0}; // @[EEPROM.scala 195:28]
  wire [2:0] _GEN_56 = done ? 3'h0 : stateReg; // @[EEPROM.scala 197:{20,31} 95:12]
  wire [16:0] _GEN_57 = sckRising ? _dataReg_T_1 : {{1'd0}, dataReg}; // @[EEPROM.scala 194:23 195:17 70:20]
  wire  _GEN_58 = sckRising ? dataReg[15] : serialReg; // @[EEPROM.scala 194:23 196:19 72:26]
  wire [2:0] _GEN_59 = sckRising ? _GEN_56 : stateReg; // @[EEPROM.scala 194:23 95:12]
  wire [16:0] _GEN_60 = 3'h7 == stateReg ? _GEN_57 : {{1'd0}, dataReg}; // @[EEPROM.scala 70:20 98:20]
  wire  _GEN_61 = 3'h7 == stateReg ? _GEN_58 : serialReg; // @[EEPROM.scala 98:20 72:26]
  wire [2:0] _GEN_62 = 3'h7 == stateReg ? _GEN_59 : stateReg; // @[EEPROM.scala 95:12 98:20]
  wire  _GEN_63 = 3'h6 == stateReg ? _GEN_53 : _GEN_61; // @[EEPROM.scala 98:20]
  wire [16:0] _GEN_64 = 3'h6 == stateReg ? _GEN_54 : _GEN_60; // @[EEPROM.scala 98:20]
  wire [2:0] _GEN_65 = 3'h6 == stateReg ? _GEN_55 : _GEN_62; // @[EEPROM.scala 98:20]
  wire [5:0] _GEN_66 = 3'h5 == stateReg ? _GEN_50 : addrReg; // @[EEPROM.scala 69:20 98:20]
  wire [2:0] _GEN_67 = 3'h5 == stateReg ? _GEN_51 : _GEN_65; // @[EEPROM.scala 98:20]
  wire  _GEN_68 = 3'h5 == stateReg ? serialReg : _GEN_63; // @[EEPROM.scala 98:20 72:26]
  wire [16:0] _GEN_69 = 3'h5 == stateReg ? {{1'd0}, dataReg} : _GEN_64; // @[EEPROM.scala 70:20 98:20]
  wire [16:0] _GEN_70 = 3'h4 == stateReg ? {{1'd0}, _GEN_46} : _GEN_69; // @[EEPROM.scala 98:20]
  wire [2:0] _GEN_71 = 3'h4 == stateReg ? _GEN_48 : _GEN_67; // @[EEPROM.scala 98:20]
  wire [5:0] _GEN_72 = 3'h4 == stateReg ? addrReg : _GEN_66; // @[EEPROM.scala 69:20 98:20]
  wire  _GEN_73 = 3'h4 == stateReg ? serialReg : _GEN_68; // @[EEPROM.scala 98:20 72:26]
  wire [16:0] _GEN_74 = 3'h3 == stateReg ? {{1'd0}, _GEN_46} : _GEN_70; // @[EEPROM.scala 98:20]
  wire [2:0] _GEN_75 = 3'h3 == stateReg ? _GEN_47 : _GEN_71; // @[EEPROM.scala 98:20]
  wire  _GEN_77 = 3'h3 == stateReg ? serialReg : _GEN_73; // @[EEPROM.scala 98:20 72:26]
  wire  _GEN_81 = 3'h2 == stateReg ? _GEN_41 : _GEN_77; // @[EEPROM.scala 98:20]
  wire [2:0] _GEN_82 = 3'h2 == stateReg ? _GEN_42 : _GEN_75; // @[EEPROM.scala 98:20]
  wire [16:0] _GEN_85 = 3'h2 == stateReg ? {{1'd0}, dataReg} : _GEN_74; // @[EEPROM.scala 70:20 98:20]
  wire  _GEN_90 = 3'h1 == stateReg ? serialReg : _GEN_81; // @[EEPROM.scala 98:20 72:26]
  wire [16:0] _GEN_93 = 3'h1 == stateReg ? {{1'd0}, dataReg} : _GEN_85; // @[EEPROM.scala 70:20 98:20]
  wire [16:0] _GEN_96 = 3'h0 == stateReg ? 17'hffff : _GEN_93; // @[EEPROM.scala 103:15 98:20]
  wire  _GEN_97 = 3'h0 == stateReg | _GEN_90; // @[EEPROM.scala 104:17 98:20]
  assign io_mem_rd = stateReg == 3'h3; // @[EEPROM.scala 207:25]
  assign io_mem_wr = stateReg == 3'h5; // @[EEPROM.scala 208:25]
  assign io_mem_addr = {addrReg,1'h0}; // @[EEPROM.scala 209:26]
  assign io_mem_din = dataReg; // @[EEPROM.scala 211:14]
  assign io_serial_sdo = serialReg; // @[EEPROM.scala 206:17]
  always @(posedge clock) begin
    if (reset) begin // @[EEPROM.scala 65:25]
      stateReg <= 3'h0; // @[EEPROM.scala 65:25]
    end else if (~io_serial_cs) begin // @[EEPROM.scala 203:23]
      stateReg <= 3'h0; // @[EEPROM.scala 203:34]
    end else if (3'h0 == stateReg) begin // @[EEPROM.scala 98:20]
      if (io_serial_cs) begin // @[EEPROM.scala 106:26]
        stateReg <= 3'h1; // @[EEPROM.scala 106:37]
      end
    end else if (3'h1 == stateReg) begin // @[EEPROM.scala 98:20]
      stateReg <= _GEN_2;
    end else begin
      stateReg <= _GEN_82;
    end
    if (reset) begin // @[EEPROM.scala 68:27]
      counterReg <= 17'h0; // @[EEPROM.scala 68:27]
    end else if (3'h0 == stateReg) begin // @[EEPROM.scala 98:20]
      counterReg <= 17'h80; // @[EEPROM.scala 101:18]
    end else if (3'h1 == stateReg) begin // @[EEPROM.scala 98:20]
      counterReg <= _GEN_0;
    end else if (3'h2 == stateReg) begin // @[EEPROM.scala 98:20]
      counterReg <= _GEN_40;
    end else begin
      counterReg <= _GEN_0;
    end
    if (3'h0 == stateReg) begin // @[EEPROM.scala 98:20]
      addrReg <= 6'h0; // @[EEPROM.scala 102:15]
    end else if (!(3'h1 == stateReg)) begin // @[EEPROM.scala 98:20]
      if (3'h2 == stateReg) begin // @[EEPROM.scala 98:20]
        if (sckRising) begin // @[EEPROM.scala 116:23]
          addrReg <= _GEN_35;
        end
      end else if (!(3'h3 == stateReg)) begin // @[EEPROM.scala 98:20]
        addrReg <= _GEN_72;
      end
    end
    dataReg <= _GEN_96[15:0];
    if (!(3'h0 == stateReg)) begin // @[EEPROM.scala 98:20]
      if (!(3'h1 == stateReg)) begin // @[EEPROM.scala 98:20]
        if (3'h2 == stateReg) begin // @[EEPROM.scala 98:20]
          if (sckRising) begin // @[EEPROM.scala 116:23]
            opcodeReg <= data[6:5]; // @[EEPROM.scala 120:19]
          end
        end
      end
    end
    serialReg <= reset | _GEN_97; // @[EEPROM.scala 72:{26,26}]
    if (reset) begin // @[EEPROM.scala 73:28]
      writeAllReg <= 1'h0; // @[EEPROM.scala 73:28]
    end else if (3'h0 == stateReg) begin // @[EEPROM.scala 98:20]
      writeAllReg <= 1'h0; // @[EEPROM.scala 105:19]
    end else if (!(3'h1 == stateReg)) begin // @[EEPROM.scala 98:20]
      if (3'h2 == stateReg) begin // @[EEPROM.scala 98:20]
        writeAllReg <= _GEN_43;
      end
    end
    if (reset) begin // @[EEPROM.scala 74:31]
      writeEnableReg <= 1'h0; // @[EEPROM.scala 74:31]
    end else if (!(3'h0 == stateReg)) begin // @[EEPROM.scala 98:20]
      if (!(3'h1 == stateReg)) begin // @[EEPROM.scala 98:20]
        if (3'h2 == stateReg) begin // @[EEPROM.scala 98:20]
          writeEnableReg <= _GEN_44;
        end
      end
    end
    sckRising_REG <= io_serial_sck; // @[Util.scala 158:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  counterReg = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  addrReg = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  dataReg = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  opcodeReg = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  serialReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  writeAllReg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  writeEnableReg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sckRising_REG = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SinglePortRam(
  input         clock,
  input         io_rd,
  input         io_wr,
  input  [14:0] io_addr,
  input  [1:0]  io_mask,
  input  [15:0] io_din,
  output [15:0] io_dout
);
  wire  ram_clk; // @[SinglePortRam.scala 72:19]
  wire  ram_rd; // @[SinglePortRam.scala 72:19]
  wire  ram_wr; // @[SinglePortRam.scala 72:19]
  wire [14:0] ram_addr; // @[SinglePortRam.scala 72:19]
  wire [1:0] ram_mask; // @[SinglePortRam.scala 72:19]
  wire [15:0] ram_din; // @[SinglePortRam.scala 72:19]
  wire [15:0] ram_dout; // @[SinglePortRam.scala 72:19]
  single_port_ram #(.ADDR_WIDTH(15), .DATA_WIDTH(16), .DEPTH(0), .MASK_ENABLE("TRUE")) ram ( // @[SinglePortRam.scala 72:19]
    .clk(ram_clk),
    .rd(ram_rd),
    .wr(ram_wr),
    .addr(ram_addr),
    .mask(ram_mask),
    .din(ram_din),
    .dout(ram_dout)
  );
  assign io_dout = ram_dout; // @[SinglePortRam.scala 79:11]
  assign ram_clk = clock; // @[SinglePortRam.scala 73:14]
  assign ram_rd = io_rd; // @[SinglePortRam.scala 74:13]
  assign ram_wr = io_wr; // @[SinglePortRam.scala 75:13]
  assign ram_addr = io_addr; // @[SinglePortRam.scala 76:15]
  assign ram_mask = io_mask; // @[SinglePortRam.scala 77:15]
  assign ram_din = io_din; // @[SinglePortRam.scala 78:14]
endmodule
module TrueDualPortRam(
  input          clock,
  input          io_clockB,
  input          io_portA_rd,
  input          io_portA_wr,
  input  [14:0]  io_portA_addr,
  input  [1:0]   io_portA_mask,
  input  [15:0]  io_portA_din,
  output [15:0]  io_portA_dout,
  input          io_portB_rd,
  input  [11:0]  io_portB_addr,
  output [127:0] io_portB_dout
);
  wire  ram_clk_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_rd_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_wr_a; // @[TrueDualPortRam.scala 99:19]
  wire [14:0] ram_addr_a; // @[TrueDualPortRam.scala 99:19]
  wire [1:0] ram_mask_a; // @[TrueDualPortRam.scala 99:19]
  wire [15:0] ram_din_a; // @[TrueDualPortRam.scala 99:19]
  wire [15:0] ram_dout_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_clk_b; // @[TrueDualPortRam.scala 99:19]
  wire  ram_rd_b; // @[TrueDualPortRam.scala 99:19]
  wire [11:0] ram_addr_b; // @[TrueDualPortRam.scala 99:19]
  wire [127:0] ram_dout_b; // @[TrueDualPortRam.scala 99:19]
  true_dual_port_ram
    #(.ADDR_WIDTH_A(15), .DEPTH_B(0), .DEPTH_A(0), .DATA_WIDTH_A(16), .DATA_WIDTH_B(128), .MASK_ENABLE("TRUE"), .ADDR_WIDTH_B(12))
    ram ( // @[TrueDualPortRam.scala 99:19]
    .clk_a(ram_clk_a),
    .rd_a(ram_rd_a),
    .wr_a(ram_wr_a),
    .addr_a(ram_addr_a),
    .mask_a(ram_mask_a),
    .din_a(ram_din_a),
    .dout_a(ram_dout_a),
    .clk_b(ram_clk_b),
    .rd_b(ram_rd_b),
    .addr_b(ram_addr_b),
    .dout_b(ram_dout_b)
  );
  assign io_portA_dout = ram_dout_a; // @[TrueDualPortRam.scala 106:17]
  assign io_portB_dout = ram_dout_b; // @[TrueDualPortRam.scala 110:17]
  assign ram_clk_a = clock; // @[TrueDualPortRam.scala 100:16]
  assign ram_rd_a = io_portA_rd; // @[TrueDualPortRam.scala 101:15]
  assign ram_wr_a = io_portA_wr; // @[TrueDualPortRam.scala 102:15]
  assign ram_addr_a = io_portA_addr; // @[TrueDualPortRam.scala 103:17]
  assign ram_mask_a = io_portA_mask; // @[TrueDualPortRam.scala 104:17]
  assign ram_din_a = io_portA_din; // @[TrueDualPortRam.scala 105:16]
  assign ram_clk_b = io_clockB; // @[TrueDualPortRam.scala 107:16]
  assign ram_rd_b = io_portB_rd; // @[TrueDualPortRam.scala 108:15]
  assign ram_addr_b = io_portB_addr; // @[TrueDualPortRam.scala 109:17]
endmodule
module TrueDualPortRam_1(
  input         clock,
  input         io_clockB,
  input         io_portA_rd,
  input         io_portA_wr,
  input  [12:0] io_portA_addr,
  input  [1:0]  io_portA_mask,
  input  [15:0] io_portA_din,
  output [15:0] io_portA_dout,
  input  [11:0] io_portB_addr,
  output [31:0] io_portB_dout
);
  wire  ram_clk_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_rd_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_wr_a; // @[TrueDualPortRam.scala 99:19]
  wire [12:0] ram_addr_a; // @[TrueDualPortRam.scala 99:19]
  wire [1:0] ram_mask_a; // @[TrueDualPortRam.scala 99:19]
  wire [15:0] ram_din_a; // @[TrueDualPortRam.scala 99:19]
  wire [15:0] ram_dout_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_clk_b; // @[TrueDualPortRam.scala 99:19]
  wire  ram_rd_b; // @[TrueDualPortRam.scala 99:19]
  wire [11:0] ram_addr_b; // @[TrueDualPortRam.scala 99:19]
  wire [31:0] ram_dout_b; // @[TrueDualPortRam.scala 99:19]
  true_dual_port_ram
    #(.ADDR_WIDTH_A(13), .DEPTH_B(0), .DEPTH_A(0), .DATA_WIDTH_A(16), .DATA_WIDTH_B(32), .MASK_ENABLE("TRUE"), .ADDR_WIDTH_B(12))
    ram ( // @[TrueDualPortRam.scala 99:19]
    .clk_a(ram_clk_a),
    .rd_a(ram_rd_a),
    .wr_a(ram_wr_a),
    .addr_a(ram_addr_a),
    .mask_a(ram_mask_a),
    .din_a(ram_din_a),
    .dout_a(ram_dout_a),
    .clk_b(ram_clk_b),
    .rd_b(ram_rd_b),
    .addr_b(ram_addr_b),
    .dout_b(ram_dout_b)
  );
  assign io_portA_dout = ram_dout_a; // @[TrueDualPortRam.scala 106:17]
  assign io_portB_dout = ram_dout_b; // @[TrueDualPortRam.scala 110:17]
  assign ram_clk_a = clock; // @[TrueDualPortRam.scala 100:16]
  assign ram_rd_a = io_portA_rd; // @[TrueDualPortRam.scala 101:15]
  assign ram_wr_a = io_portA_wr; // @[TrueDualPortRam.scala 102:15]
  assign ram_addr_a = io_portA_addr; // @[TrueDualPortRam.scala 103:17]
  assign ram_mask_a = io_portA_mask; // @[TrueDualPortRam.scala 104:17]
  assign ram_din_a = io_portA_din; // @[TrueDualPortRam.scala 105:16]
  assign ram_clk_b = io_clockB; // @[TrueDualPortRam.scala 107:16]
  assign ram_rd_b = 1'h1; // @[TrueDualPortRam.scala 108:15]
  assign ram_addr_b = io_portB_addr; // @[TrueDualPortRam.scala 109:17]
endmodule
module TrueDualPortRam_4(
  input         clock,
  input         io_clockB,
  input         io_portA_rd,
  input         io_portA_wr,
  input  [10:0] io_portA_addr,
  input  [1:0]  io_portA_mask,
  input  [15:0] io_portA_din,
  output [15:0] io_portA_dout,
  input  [9:0]  io_portB_addr,
  output [31:0] io_portB_dout
);
  wire  ram_clk_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_rd_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_wr_a; // @[TrueDualPortRam.scala 99:19]
  wire [10:0] ram_addr_a; // @[TrueDualPortRam.scala 99:19]
  wire [1:0] ram_mask_a; // @[TrueDualPortRam.scala 99:19]
  wire [15:0] ram_din_a; // @[TrueDualPortRam.scala 99:19]
  wire [15:0] ram_dout_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_clk_b; // @[TrueDualPortRam.scala 99:19]
  wire  ram_rd_b; // @[TrueDualPortRam.scala 99:19]
  wire [9:0] ram_addr_b; // @[TrueDualPortRam.scala 99:19]
  wire [31:0] ram_dout_b; // @[TrueDualPortRam.scala 99:19]
  true_dual_port_ram
    #(.ADDR_WIDTH_A(11), .DEPTH_B(0), .DEPTH_A(0), .DATA_WIDTH_A(16), .DATA_WIDTH_B(32), .MASK_ENABLE("TRUE"), .ADDR_WIDTH_B(10))
    ram ( // @[TrueDualPortRam.scala 99:19]
    .clk_a(ram_clk_a),
    .rd_a(ram_rd_a),
    .wr_a(ram_wr_a),
    .addr_a(ram_addr_a),
    .mask_a(ram_mask_a),
    .din_a(ram_din_a),
    .dout_a(ram_dout_a),
    .clk_b(ram_clk_b),
    .rd_b(ram_rd_b),
    .addr_b(ram_addr_b),
    .dout_b(ram_dout_b)
  );
  assign io_portA_dout = ram_dout_a; // @[TrueDualPortRam.scala 106:17]
  assign io_portB_dout = ram_dout_b; // @[TrueDualPortRam.scala 110:17]
  assign ram_clk_a = clock; // @[TrueDualPortRam.scala 100:16]
  assign ram_rd_a = io_portA_rd; // @[TrueDualPortRam.scala 101:15]
  assign ram_wr_a = io_portA_wr; // @[TrueDualPortRam.scala 102:15]
  assign ram_addr_a = io_portA_addr; // @[TrueDualPortRam.scala 103:17]
  assign ram_mask_a = io_portA_mask; // @[TrueDualPortRam.scala 104:17]
  assign ram_din_a = io_portA_din; // @[TrueDualPortRam.scala 105:16]
  assign ram_clk_b = io_clockB; // @[TrueDualPortRam.scala 107:16]
  assign ram_rd_b = 1'h1; // @[TrueDualPortRam.scala 108:15]
  assign ram_addr_b = io_portB_addr; // @[TrueDualPortRam.scala 109:17]
endmodule
module TrueDualPortRam_7(
  input         clock,
  input         io_clockB,
  input         io_portA_rd,
  input         io_portA_wr,
  input  [9:0]  io_portA_addr,
  input  [1:0]  io_portA_mask,
  input  [15:0] io_portA_din,
  output [15:0] io_portA_dout,
  input  [8:0]  io_portB_addr,
  output [31:0] io_portB_dout
);
  wire  ram_clk_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_rd_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_wr_a; // @[TrueDualPortRam.scala 99:19]
  wire [9:0] ram_addr_a; // @[TrueDualPortRam.scala 99:19]
  wire [1:0] ram_mask_a; // @[TrueDualPortRam.scala 99:19]
  wire [15:0] ram_din_a; // @[TrueDualPortRam.scala 99:19]
  wire [15:0] ram_dout_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_clk_b; // @[TrueDualPortRam.scala 99:19]
  wire  ram_rd_b; // @[TrueDualPortRam.scala 99:19]
  wire [8:0] ram_addr_b; // @[TrueDualPortRam.scala 99:19]
  wire [31:0] ram_dout_b; // @[TrueDualPortRam.scala 99:19]
  true_dual_port_ram
    #(.ADDR_WIDTH_A(10), .DEPTH_B(0), .DEPTH_A(0), .DATA_WIDTH_A(16), .DATA_WIDTH_B(32), .MASK_ENABLE("TRUE"), .ADDR_WIDTH_B(9))
    ram ( // @[TrueDualPortRam.scala 99:19]
    .clk_a(ram_clk_a),
    .rd_a(ram_rd_a),
    .wr_a(ram_wr_a),
    .addr_a(ram_addr_a),
    .mask_a(ram_mask_a),
    .din_a(ram_din_a),
    .dout_a(ram_dout_a),
    .clk_b(ram_clk_b),
    .rd_b(ram_rd_b),
    .addr_b(ram_addr_b),
    .dout_b(ram_dout_b)
  );
  assign io_portA_dout = ram_dout_a; // @[TrueDualPortRam.scala 106:17]
  assign io_portB_dout = ram_dout_b; // @[TrueDualPortRam.scala 110:17]
  assign ram_clk_a = clock; // @[TrueDualPortRam.scala 100:16]
  assign ram_rd_a = io_portA_rd; // @[TrueDualPortRam.scala 101:15]
  assign ram_wr_a = io_portA_wr; // @[TrueDualPortRam.scala 102:15]
  assign ram_addr_a = io_portA_addr; // @[TrueDualPortRam.scala 103:17]
  assign ram_mask_a = io_portA_mask; // @[TrueDualPortRam.scala 104:17]
  assign ram_din_a = io_portA_din; // @[TrueDualPortRam.scala 105:16]
  assign ram_clk_b = io_clockB; // @[TrueDualPortRam.scala 107:16]
  assign ram_rd_b = 1'h1; // @[TrueDualPortRam.scala 108:15]
  assign ram_addr_b = io_portB_addr; // @[TrueDualPortRam.scala 109:17]
endmodule
module TrueDualPortRam_10(
  input         clock,
  input         io_clockB,
  input         io_portA_rd,
  input         io_portA_wr,
  input  [14:0] io_portA_addr,
  input  [1:0]  io_portA_mask,
  input  [15:0] io_portA_din,
  output [15:0] io_portA_dout,
  input  [14:0] io_portB_addr,
  output [15:0] io_portB_dout
);
  wire  ram_clk_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_rd_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_wr_a; // @[TrueDualPortRam.scala 99:19]
  wire [14:0] ram_addr_a; // @[TrueDualPortRam.scala 99:19]
  wire [1:0] ram_mask_a; // @[TrueDualPortRam.scala 99:19]
  wire [15:0] ram_din_a; // @[TrueDualPortRam.scala 99:19]
  wire [15:0] ram_dout_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_clk_b; // @[TrueDualPortRam.scala 99:19]
  wire  ram_rd_b; // @[TrueDualPortRam.scala 99:19]
  wire [14:0] ram_addr_b; // @[TrueDualPortRam.scala 99:19]
  wire [15:0] ram_dout_b; // @[TrueDualPortRam.scala 99:19]
  true_dual_port_ram
    #(.ADDR_WIDTH_A(15), .DEPTH_B(0), .DEPTH_A(0), .DATA_WIDTH_A(16), .DATA_WIDTH_B(16), .MASK_ENABLE("TRUE"), .ADDR_WIDTH_B(15))
    ram ( // @[TrueDualPortRam.scala 99:19]
    .clk_a(ram_clk_a),
    .rd_a(ram_rd_a),
    .wr_a(ram_wr_a),
    .addr_a(ram_addr_a),
    .mask_a(ram_mask_a),
    .din_a(ram_din_a),
    .dout_a(ram_dout_a),
    .clk_b(ram_clk_b),
    .rd_b(ram_rd_b),
    .addr_b(ram_addr_b),
    .dout_b(ram_dout_b)
  );
  assign io_portA_dout = ram_dout_a; // @[TrueDualPortRam.scala 106:17]
  assign io_portB_dout = ram_dout_b; // @[TrueDualPortRam.scala 110:17]
  assign ram_clk_a = clock; // @[TrueDualPortRam.scala 100:16]
  assign ram_rd_a = io_portA_rd; // @[TrueDualPortRam.scala 101:15]
  assign ram_wr_a = io_portA_wr; // @[TrueDualPortRam.scala 102:15]
  assign ram_addr_a = io_portA_addr; // @[TrueDualPortRam.scala 103:17]
  assign ram_mask_a = io_portA_mask; // @[TrueDualPortRam.scala 104:17]
  assign ram_din_a = io_portA_din; // @[TrueDualPortRam.scala 105:16]
  assign ram_clk_b = io_clockB; // @[TrueDualPortRam.scala 107:16]
  assign ram_rd_b = 1'h1; // @[TrueDualPortRam.scala 108:15]
  assign ram_addr_b = io_portB_addr; // @[TrueDualPortRam.scala 109:17]
endmodule
module RegisterFile_2(
  input         clock,
  input         io_mem_wr,
  input  [1:0]  io_mem_addr,
  input  [1:0]  io_mem_mask,
  input  [15:0] io_mem_din,
  output [15:0] io_mem_dout,
  output [15:0] io_regs_0,
  output [15:0] io_regs_1,
  output [15:0] io_regs_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] regs_0; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_1; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_2; // @[RegisterFile.scala 56:17]
  wire [15:0] _GEN_1 = 2'h1 == io_mem_addr ? regs_1 : regs_0; // @[]
  wire [15:0] _GEN_2 = 2'h2 == io_mem_addr ? regs_2 : _GEN_1; // @[]
  wire [7:0] bytes_0 = io_mem_wr & io_mem_mask[0] ? io_mem_din[7:0] : _GEN_2[7:0]; // @[RegisterFile.scala 62:28 66:{39,50}]
  wire [7:0] bytes_1 = io_mem_wr & io_mem_mask[1] ? io_mem_din[15:8] : _GEN_2[15:8]; // @[RegisterFile.scala 62:28 66:{39,50}]
  wire [15:0] _regs_T = {bytes_1,bytes_0}; // @[RegisterFile.scala 70:17]
  assign io_mem_dout = 2'h2 == io_mem_addr ? regs_2 : _GEN_1; // @[]
  assign io_regs_0 = regs_0; // @[RegisterFile.scala 74:11]
  assign io_regs_1 = regs_1; // @[RegisterFile.scala 74:11]
  assign io_regs_2 = regs_2; // @[RegisterFile.scala 74:11]
  always @(posedge clock) begin
    if (2'h0 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_0 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (2'h1 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_1 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (2'h2 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_2 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegisterFile_5(
  input         clock,
  input         io_mem_wr,
  input  [2:0]  io_mem_addr,
  input  [1:0]  io_mem_mask,
  input  [15:0] io_mem_din,
  output [15:0] io_regs_0,
  output [15:0] io_regs_1,
  output [15:0] io_regs_4,
  output [15:0] io_regs_5
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] regs_0; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_1; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_2; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_3; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_4; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_5; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_6; // @[RegisterFile.scala 56:17]
  reg [15:0] regs_7; // @[RegisterFile.scala 56:17]
  wire [15:0] _GEN_1 = 3'h1 == io_mem_addr ? regs_1 : regs_0; // @[]
  wire [15:0] _GEN_2 = 3'h2 == io_mem_addr ? regs_2 : _GEN_1; // @[]
  wire [15:0] _GEN_3 = 3'h3 == io_mem_addr ? regs_3 : _GEN_2; // @[]
  wire [15:0] _GEN_4 = 3'h4 == io_mem_addr ? regs_4 : _GEN_3; // @[]
  wire [15:0] _GEN_5 = 3'h5 == io_mem_addr ? regs_5 : _GEN_4; // @[]
  wire [15:0] _GEN_6 = 3'h6 == io_mem_addr ? regs_6 : _GEN_5; // @[]
  wire [15:0] _GEN_7 = 3'h7 == io_mem_addr ? regs_7 : _GEN_6; // @[]
  wire [7:0] bytes_0 = io_mem_wr & io_mem_mask[0] ? io_mem_din[7:0] : _GEN_7[7:0]; // @[RegisterFile.scala 62:28 66:{39,50}]
  wire [7:0] bytes_1 = io_mem_wr & io_mem_mask[1] ? io_mem_din[15:8] : _GEN_7[15:8]; // @[RegisterFile.scala 62:28 66:{39,50}]
  wire [15:0] _regs_T = {bytes_1,bytes_0}; // @[RegisterFile.scala 70:17]
  assign io_regs_0 = regs_0; // @[RegisterFile.scala 74:11]
  assign io_regs_1 = regs_1; // @[RegisterFile.scala 74:11]
  assign io_regs_4 = regs_4; // @[RegisterFile.scala 74:11]
  assign io_regs_5 = regs_5; // @[RegisterFile.scala 74:11]
  always @(posedge clock) begin
    if (3'h0 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_0 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h1 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_1 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h2 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_2 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h3 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_3 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h4 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_4 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h5 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_5 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h6 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_6 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
    if (3'h7 == io_mem_addr) begin // @[RegisterFile.scala 70:8]
      regs_7 <= _regs_T; // @[RegisterFile.scala 70:8]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Main(
  input          clock,
  input          reset,
  input          io_videoClock,
  input          io_spriteClock,
  input  [3:0]   io_gameIndex,
  input          io_options_service,
  input          io_player_0_up,
  input          io_player_0_down,
  input          io_player_0_left,
  input          io_player_0_right,
  input  [3:0]   io_player_0_buttons,
  input          io_player_0_start,
  input          io_player_0_coin,
  input          io_player_0_pause,
  input          io_player_1_up,
  input          io_player_1_down,
  input          io_player_1_left,
  input          io_player_1_right,
  input  [3:0]   io_player_1_buttons,
  input          io_player_1_start,
  input          io_player_1_coin,
  input          io_player_1_pause,
  input  [15:0]  io_dips_0,
  input          io_video_vBlank,
  output         io_gpuMem_layer_0_regs_tileSize,
  output         io_gpuMem_layer_0_regs_enable,
  output         io_gpuMem_layer_0_regs_flipX,
  output         io_gpuMem_layer_0_regs_flipY,
  output         io_gpuMem_layer_0_regs_rowScrollEnable,
  output         io_gpuMem_layer_0_regs_rowSelectEnable,
  output [8:0]   io_gpuMem_layer_0_regs_scroll_x,
  output [8:0]   io_gpuMem_layer_0_regs_scroll_y,
  input  [11:0]  io_gpuMem_layer_0_vram8x8_addr,
  output [31:0]  io_gpuMem_layer_0_vram8x8_dout,
  input  [9:0]   io_gpuMem_layer_0_vram16x16_addr,
  output [31:0]  io_gpuMem_layer_0_vram16x16_dout,
  input  [8:0]   io_gpuMem_layer_0_lineRam_addr,
  output [31:0]  io_gpuMem_layer_0_lineRam_dout,
  output         io_gpuMem_layer_1_regs_tileSize,
  output         io_gpuMem_layer_1_regs_enable,
  output         io_gpuMem_layer_1_regs_flipX,
  output         io_gpuMem_layer_1_regs_flipY,
  output         io_gpuMem_layer_1_regs_rowScrollEnable,
  output         io_gpuMem_layer_1_regs_rowSelectEnable,
  output [8:0]   io_gpuMem_layer_1_regs_scroll_x,
  output [8:0]   io_gpuMem_layer_1_regs_scroll_y,
  input  [11:0]  io_gpuMem_layer_1_vram8x8_addr,
  output [31:0]  io_gpuMem_layer_1_vram8x8_dout,
  input  [9:0]   io_gpuMem_layer_1_vram16x16_addr,
  output [31:0]  io_gpuMem_layer_1_vram16x16_dout,
  input  [8:0]   io_gpuMem_layer_1_lineRam_addr,
  output [31:0]  io_gpuMem_layer_1_lineRam_dout,
  output         io_gpuMem_layer_2_regs_tileSize,
  output         io_gpuMem_layer_2_regs_enable,
  output         io_gpuMem_layer_2_regs_flipX,
  output         io_gpuMem_layer_2_regs_flipY,
  output         io_gpuMem_layer_2_regs_rowScrollEnable,
  output         io_gpuMem_layer_2_regs_rowSelectEnable,
  output [8:0]   io_gpuMem_layer_2_regs_scroll_x,
  output [8:0]   io_gpuMem_layer_2_regs_scroll_y,
  input  [11:0]  io_gpuMem_layer_2_vram8x8_addr,
  output [31:0]  io_gpuMem_layer_2_vram8x8_dout,
  input  [9:0]   io_gpuMem_layer_2_vram16x16_addr,
  output [31:0]  io_gpuMem_layer_2_vram16x16_dout,
  input  [8:0]   io_gpuMem_layer_2_lineRam_addr,
  output [31:0]  io_gpuMem_layer_2_lineRam_dout,
  output [8:0]   io_gpuMem_sprite_regs_offset_x,
  output [8:0]   io_gpuMem_sprite_regs_offset_y,
  output [1:0]   io_gpuMem_sprite_regs_bank,
  output         io_gpuMem_sprite_regs_fixed,
  output         io_gpuMem_sprite_regs_hFlip,
  input          io_gpuMem_sprite_vram_rd,
  input  [11:0]  io_gpuMem_sprite_vram_addr,
  output [127:0] io_gpuMem_sprite_vram_dout,
  input  [14:0]  io_gpuMem_paletteRam_addr,
  output [15:0]  io_gpuMem_paletteRam_dout,
  output         io_soundCtrl_oki_0_wr,
  output [15:0]  io_soundCtrl_oki_0_din,
  input  [15:0]  io_soundCtrl_oki_0_dout,
  output         io_soundCtrl_oki_1_wr,
  output [15:0]  io_soundCtrl_oki_1_din,
  input  [15:0]  io_soundCtrl_oki_1_dout,
  output         io_soundCtrl_nmk_wr,
  output [22:0]  io_soundCtrl_nmk_addr,
  output [15:0]  io_soundCtrl_nmk_din,
  output         io_soundCtrl_ymz_rd,
  output         io_soundCtrl_ymz_wr,
  output [22:0]  io_soundCtrl_ymz_addr,
  output [15:0]  io_soundCtrl_ymz_din,
  input  [15:0]  io_soundCtrl_ymz_dout,
  output         io_soundCtrl_req,
  output [15:0]  io_soundCtrl_data,
  input          io_soundCtrl_irq,
  output         io_progRom_rd,
  output [19:0]  io_progRom_addr,
  input  [15:0]  io_progRom_dout,
  input          io_progRom_valid,
  output         io_eeprom_rd,
  output         io_eeprom_wr,
  output [6:0]   io_eeprom_addr,
  output [15:0]  io_eeprom_din,
  input  [15:0]  io_eeprom_dout,
  input          io_eeprom_wait_n,
  input          io_eeprom_valid,
  output         io_spriteFrameBufferSwap
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
`endif // RANDOMIZE_REG_INIT
  wire  cpu_clock; // @[Main.scala 91:19]
  wire  cpu_reset; // @[Main.scala 91:19]
  wire  cpu_io_halt; // @[Main.scala 91:19]
  wire  cpu_io_as; // @[Main.scala 91:19]
  wire  cpu_io_rw; // @[Main.scala 91:19]
  wire  cpu_io_uds; // @[Main.scala 91:19]
  wire  cpu_io_lds; // @[Main.scala 91:19]
  wire  cpu_io_dtack; // @[Main.scala 91:19]
  wire  cpu_io_vpa; // @[Main.scala 91:19]
  wire [2:0] cpu_io_ipl; // @[Main.scala 91:19]
  wire [2:0] cpu_io_fc; // @[Main.scala 91:19]
  wire [22:0] cpu_io_addr; // @[Main.scala 91:19]
  wire [15:0] cpu_io_din; // @[Main.scala 91:19]
  wire [15:0] cpu_io_dout; // @[Main.scala 91:19]
  wire  eeprom_clock; // @[Main.scala 109:22]
  wire  eeprom_reset; // @[Main.scala 109:22]
  wire  eeprom_io_mem_rd; // @[Main.scala 109:22]
  wire  eeprom_io_mem_wr; // @[Main.scala 109:22]
  wire [6:0] eeprom_io_mem_addr; // @[Main.scala 109:22]
  wire [15:0] eeprom_io_mem_din; // @[Main.scala 109:22]
  wire [15:0] eeprom_io_mem_dout; // @[Main.scala 109:22]
  wire  eeprom_io_mem_wait_n; // @[Main.scala 109:22]
  wire  eeprom_io_mem_valid; // @[Main.scala 109:22]
  wire  eeprom_io_serial_cs; // @[Main.scala 109:22]
  wire  eeprom_io_serial_sck; // @[Main.scala 109:22]
  wire  eeprom_io_serial_sdi; // @[Main.scala 109:22]
  wire  eeprom_io_serial_sdo; // @[Main.scala 109:22]
  wire  mainRam_clock; // @[Main.scala 120:23]
  wire  mainRam_io_rd; // @[Main.scala 120:23]
  wire  mainRam_io_wr; // @[Main.scala 120:23]
  wire [14:0] mainRam_io_addr; // @[Main.scala 120:23]
  wire [1:0] mainRam_io_mask; // @[Main.scala 120:23]
  wire [15:0] mainRam_io_din; // @[Main.scala 120:23]
  wire [15:0] mainRam_io_dout; // @[Main.scala 120:23]
  wire  spriteRam_clock; // @[Main.scala 128:25]
  wire  spriteRam_io_clockB; // @[Main.scala 128:25]
  wire  spriteRam_io_portA_rd; // @[Main.scala 128:25]
  wire  spriteRam_io_portA_wr; // @[Main.scala 128:25]
  wire [14:0] spriteRam_io_portA_addr; // @[Main.scala 128:25]
  wire [1:0] spriteRam_io_portA_mask; // @[Main.scala 128:25]
  wire [15:0] spriteRam_io_portA_din; // @[Main.scala 128:25]
  wire [15:0] spriteRam_io_portA_dout; // @[Main.scala 128:25]
  wire  spriteRam_io_portB_rd; // @[Main.scala 128:25]
  wire [11:0] spriteRam_io_portB_addr; // @[Main.scala 128:25]
  wire [127:0] spriteRam_io_portB_dout; // @[Main.scala 128:25]
  wire  vram8x8_0_clock; // @[Main.scala 141:21]
  wire  vram8x8_0_io_clockB; // @[Main.scala 141:21]
  wire  vram8x8_0_io_portA_rd; // @[Main.scala 141:21]
  wire  vram8x8_0_io_portA_wr; // @[Main.scala 141:21]
  wire [12:0] vram8x8_0_io_portA_addr; // @[Main.scala 141:21]
  wire [1:0] vram8x8_0_io_portA_mask; // @[Main.scala 141:21]
  wire [15:0] vram8x8_0_io_portA_din; // @[Main.scala 141:21]
  wire [15:0] vram8x8_0_io_portA_dout; // @[Main.scala 141:21]
  wire [11:0] vram8x8_0_io_portB_addr; // @[Main.scala 141:21]
  wire [31:0] vram8x8_0_io_portB_dout; // @[Main.scala 141:21]
  wire  vram8x8_1_clock; // @[Main.scala 141:21]
  wire  vram8x8_1_io_clockB; // @[Main.scala 141:21]
  wire  vram8x8_1_io_portA_rd; // @[Main.scala 141:21]
  wire  vram8x8_1_io_portA_wr; // @[Main.scala 141:21]
  wire [12:0] vram8x8_1_io_portA_addr; // @[Main.scala 141:21]
  wire [1:0] vram8x8_1_io_portA_mask; // @[Main.scala 141:21]
  wire [15:0] vram8x8_1_io_portA_din; // @[Main.scala 141:21]
  wire [15:0] vram8x8_1_io_portA_dout; // @[Main.scala 141:21]
  wire [11:0] vram8x8_1_io_portB_addr; // @[Main.scala 141:21]
  wire [31:0] vram8x8_1_io_portB_dout; // @[Main.scala 141:21]
  wire  vram8x8_2_clock; // @[Main.scala 141:21]
  wire  vram8x8_2_io_clockB; // @[Main.scala 141:21]
  wire  vram8x8_2_io_portA_rd; // @[Main.scala 141:21]
  wire  vram8x8_2_io_portA_wr; // @[Main.scala 141:21]
  wire [12:0] vram8x8_2_io_portA_addr; // @[Main.scala 141:21]
  wire [1:0] vram8x8_2_io_portA_mask; // @[Main.scala 141:21]
  wire [15:0] vram8x8_2_io_portA_din; // @[Main.scala 141:21]
  wire [15:0] vram8x8_2_io_portA_dout; // @[Main.scala 141:21]
  wire [11:0] vram8x8_2_io_portB_addr; // @[Main.scala 141:21]
  wire [31:0] vram8x8_2_io_portB_dout; // @[Main.scala 141:21]
  wire  vram16x16_0_clock; // @[Main.scala 156:21]
  wire  vram16x16_0_io_clockB; // @[Main.scala 156:21]
  wire  vram16x16_0_io_portA_rd; // @[Main.scala 156:21]
  wire  vram16x16_0_io_portA_wr; // @[Main.scala 156:21]
  wire [10:0] vram16x16_0_io_portA_addr; // @[Main.scala 156:21]
  wire [1:0] vram16x16_0_io_portA_mask; // @[Main.scala 156:21]
  wire [15:0] vram16x16_0_io_portA_din; // @[Main.scala 156:21]
  wire [15:0] vram16x16_0_io_portA_dout; // @[Main.scala 156:21]
  wire [9:0] vram16x16_0_io_portB_addr; // @[Main.scala 156:21]
  wire [31:0] vram16x16_0_io_portB_dout; // @[Main.scala 156:21]
  wire  vram16x16_1_clock; // @[Main.scala 156:21]
  wire  vram16x16_1_io_clockB; // @[Main.scala 156:21]
  wire  vram16x16_1_io_portA_rd; // @[Main.scala 156:21]
  wire  vram16x16_1_io_portA_wr; // @[Main.scala 156:21]
  wire [10:0] vram16x16_1_io_portA_addr; // @[Main.scala 156:21]
  wire [1:0] vram16x16_1_io_portA_mask; // @[Main.scala 156:21]
  wire [15:0] vram16x16_1_io_portA_din; // @[Main.scala 156:21]
  wire [15:0] vram16x16_1_io_portA_dout; // @[Main.scala 156:21]
  wire [9:0] vram16x16_1_io_portB_addr; // @[Main.scala 156:21]
  wire [31:0] vram16x16_1_io_portB_dout; // @[Main.scala 156:21]
  wire  vram16x16_2_clock; // @[Main.scala 156:21]
  wire  vram16x16_2_io_clockB; // @[Main.scala 156:21]
  wire  vram16x16_2_io_portA_rd; // @[Main.scala 156:21]
  wire  vram16x16_2_io_portA_wr; // @[Main.scala 156:21]
  wire [10:0] vram16x16_2_io_portA_addr; // @[Main.scala 156:21]
  wire [1:0] vram16x16_2_io_portA_mask; // @[Main.scala 156:21]
  wire [15:0] vram16x16_2_io_portA_din; // @[Main.scala 156:21]
  wire [15:0] vram16x16_2_io_portA_dout; // @[Main.scala 156:21]
  wire [9:0] vram16x16_2_io_portB_addr; // @[Main.scala 156:21]
  wire [31:0] vram16x16_2_io_portB_dout; // @[Main.scala 156:21]
  wire  lineRam_0_clock; // @[Main.scala 171:21]
  wire  lineRam_0_io_clockB; // @[Main.scala 171:21]
  wire  lineRam_0_io_portA_rd; // @[Main.scala 171:21]
  wire  lineRam_0_io_portA_wr; // @[Main.scala 171:21]
  wire [9:0] lineRam_0_io_portA_addr; // @[Main.scala 171:21]
  wire [1:0] lineRam_0_io_portA_mask; // @[Main.scala 171:21]
  wire [15:0] lineRam_0_io_portA_din; // @[Main.scala 171:21]
  wire [15:0] lineRam_0_io_portA_dout; // @[Main.scala 171:21]
  wire [8:0] lineRam_0_io_portB_addr; // @[Main.scala 171:21]
  wire [31:0] lineRam_0_io_portB_dout; // @[Main.scala 171:21]
  wire  lineRam_1_clock; // @[Main.scala 171:21]
  wire  lineRam_1_io_clockB; // @[Main.scala 171:21]
  wire  lineRam_1_io_portA_rd; // @[Main.scala 171:21]
  wire  lineRam_1_io_portA_wr; // @[Main.scala 171:21]
  wire [9:0] lineRam_1_io_portA_addr; // @[Main.scala 171:21]
  wire [1:0] lineRam_1_io_portA_mask; // @[Main.scala 171:21]
  wire [15:0] lineRam_1_io_portA_din; // @[Main.scala 171:21]
  wire [15:0] lineRam_1_io_portA_dout; // @[Main.scala 171:21]
  wire [8:0] lineRam_1_io_portB_addr; // @[Main.scala 171:21]
  wire [31:0] lineRam_1_io_portB_dout; // @[Main.scala 171:21]
  wire  lineRam_2_clock; // @[Main.scala 171:21]
  wire  lineRam_2_io_clockB; // @[Main.scala 171:21]
  wire  lineRam_2_io_portA_rd; // @[Main.scala 171:21]
  wire  lineRam_2_io_portA_wr; // @[Main.scala 171:21]
  wire [9:0] lineRam_2_io_portA_addr; // @[Main.scala 171:21]
  wire [1:0] lineRam_2_io_portA_mask; // @[Main.scala 171:21]
  wire [15:0] lineRam_2_io_portA_din; // @[Main.scala 171:21]
  wire [15:0] lineRam_2_io_portA_dout; // @[Main.scala 171:21]
  wire [8:0] lineRam_2_io_portB_addr; // @[Main.scala 171:21]
  wire [31:0] lineRam_2_io_portB_dout; // @[Main.scala 171:21]
  wire  paletteRam_clock; // @[Main.scala 185:26]
  wire  paletteRam_io_clockB; // @[Main.scala 185:26]
  wire  paletteRam_io_portA_rd; // @[Main.scala 185:26]
  wire  paletteRam_io_portA_wr; // @[Main.scala 185:26]
  wire [14:0] paletteRam_io_portA_addr; // @[Main.scala 185:26]
  wire [1:0] paletteRam_io_portA_mask; // @[Main.scala 185:26]
  wire [15:0] paletteRam_io_portA_din; // @[Main.scala 185:26]
  wire [15:0] paletteRam_io_portA_dout; // @[Main.scala 185:26]
  wire [14:0] paletteRam_io_portB_addr; // @[Main.scala 185:26]
  wire [15:0] paletteRam_io_portB_dout; // @[Main.scala 185:26]
  wire  layerRegs_0_clock; // @[Main.scala 198:22]
  wire  layerRegs_0_io_mem_wr; // @[Main.scala 198:22]
  wire [1:0] layerRegs_0_io_mem_addr; // @[Main.scala 198:22]
  wire [1:0] layerRegs_0_io_mem_mask; // @[Main.scala 198:22]
  wire [15:0] layerRegs_0_io_mem_din; // @[Main.scala 198:22]
  wire [15:0] layerRegs_0_io_mem_dout; // @[Main.scala 198:22]
  wire [15:0] layerRegs_0_io_regs_0; // @[Main.scala 198:22]
  wire [15:0] layerRegs_0_io_regs_1; // @[Main.scala 198:22]
  wire [15:0] layerRegs_0_io_regs_2; // @[Main.scala 198:22]
  wire  layerRegs_1_clock; // @[Main.scala 198:22]
  wire  layerRegs_1_io_mem_wr; // @[Main.scala 198:22]
  wire [1:0] layerRegs_1_io_mem_addr; // @[Main.scala 198:22]
  wire [1:0] layerRegs_1_io_mem_mask; // @[Main.scala 198:22]
  wire [15:0] layerRegs_1_io_mem_din; // @[Main.scala 198:22]
  wire [15:0] layerRegs_1_io_mem_dout; // @[Main.scala 198:22]
  wire [15:0] layerRegs_1_io_regs_0; // @[Main.scala 198:22]
  wire [15:0] layerRegs_1_io_regs_1; // @[Main.scala 198:22]
  wire [15:0] layerRegs_1_io_regs_2; // @[Main.scala 198:22]
  wire  layerRegs_2_clock; // @[Main.scala 198:22]
  wire  layerRegs_2_io_mem_wr; // @[Main.scala 198:22]
  wire [1:0] layerRegs_2_io_mem_addr; // @[Main.scala 198:22]
  wire [1:0] layerRegs_2_io_mem_mask; // @[Main.scala 198:22]
  wire [15:0] layerRegs_2_io_mem_din; // @[Main.scala 198:22]
  wire [15:0] layerRegs_2_io_mem_dout; // @[Main.scala 198:22]
  wire [15:0] layerRegs_2_io_regs_0; // @[Main.scala 198:22]
  wire [15:0] layerRegs_2_io_regs_1; // @[Main.scala 198:22]
  wire [15:0] layerRegs_2_io_regs_2; // @[Main.scala 198:22]
  wire  spriteRegs_clock; // @[Main.scala 205:26]
  wire  spriteRegs_io_mem_wr; // @[Main.scala 205:26]
  wire [2:0] spriteRegs_io_mem_addr; // @[Main.scala 205:26]
  wire [1:0] spriteRegs_io_mem_mask; // @[Main.scala 205:26]
  wire [15:0] spriteRegs_io_mem_din; // @[Main.scala 205:26]
  wire [15:0] spriteRegs_io_regs_0; // @[Main.scala 205:26]
  wire [15:0] spriteRegs_io_regs_1; // @[Main.scala 205:26]
  wire [15:0] spriteRegs_io_regs_4; // @[Main.scala 205:26]
  wire [15:0] spriteRegs_io_regs_5; // @[Main.scala 205:26]
  reg  vBlank_r; // @[Reg.scala 19:16]
  reg  vBlank; // @[Reg.scala 19:16]
  reg  vBlankRising_REG; // @[Util.scala 158:44]
  wire  vBlankRising = vBlank & ~vBlankRising_REG; // @[Util.scala 158:33]
  wire  _pauseReg_T = io_player_0_pause | io_player_1_pause; // @[Main.scala 83:61]
  reg  pauseReg_REG; // @[Util.scala 158:44]
  wire  _pauseReg_T_2 = _pauseReg_T & ~pauseReg_REG; // @[Util.scala 158:33]
  reg  pauseReg; // @[Util.scala 242:26]
  reg  videoIrq; // @[Main.scala 86:25]
  reg  agalletIrq; // @[Main.scala 87:27]
  reg [15:0] dinReg; // @[MemMap.scala 48:23]
  reg  dtackReg; // @[MemMap.scala 49:25]
  reg  readStrobe_REG; // @[Util.scala 158:44]
  wire  _readStrobe_T_1 = cpu_io_as & ~readStrobe_REG; // @[Util.scala 158:33]
  wire  readStrobe = _readStrobe_T_1 & cpu_io_rw; // @[MemMap.scala 52:40]
  reg  upperWriteStrobe_REG; // @[Util.scala 158:44]
  wire  _upperWriteStrobe_T_1 = cpu_io_uds & ~upperWriteStrobe_REG; // @[Util.scala 158:33]
  wire  _upperWriteStrobe_T_3 = ~cpu_io_rw; // @[MemMap.scala 53:60]
  wire  upperWriteStrobe = cpu_io_as & _upperWriteStrobe_T_1 & ~cpu_io_rw; // @[MemMap.scala 53:57]
  reg  lowerWriteStrobe_REG; // @[Util.scala 158:44]
  wire  _lowerWriteStrobe_T_1 = cpu_io_lds & ~lowerWriteStrobe_REG; // @[Util.scala 158:33]
  wire  lowerWriteStrobe = cpu_io_as & _lowerWriteStrobe_T_1 & _upperWriteStrobe_T_3; // @[MemMap.scala 54:57]
  wire  writeStrobe = upperWriteStrobe | lowerWriteStrobe; // @[MemMap.scala 55:38]
  wire  _cpu_io_ipl_T = videoIrq | io_soundCtrl_irq; // @[Main.scala 96:26]
  wire  _cs_T = io_gameIndex == 4'h5; // @[Main.scala 111:29]
  wire  _T_260 = io_gameIndex == 4'h7; // @[Main.scala 393:21]
  wire [15:0] _GEN_193 = cpu_io_dout; // @[Main.scala 267:42 MemMap.scala 107:15]
  wire [15:0] _GEN_350 = io_gameIndex == 4'h2 ? cpu_io_dout : _GEN_193; // @[Main.scala 285:42 MemMap.scala 107:15]
  wire [15:0] _GEN_518 = io_gameIndex == 4'h1 ? cpu_io_dout : _GEN_350; // @[Main.scala 306:42 MemMap.scala 107:15]
  wire [15:0] _GEN_704 = io_gameIndex == 4'h3 ? cpu_io_dout : _GEN_518; // @[Main.scala 326:41 MemMap.scala 107:15]
  wire [15:0] _GEN_1175 = _cs_T ? cpu_io_dout : _GEN_704; // @[Main.scala 368:41 MemMap.scala 153:15]
  wire [15:0] _GEN_1368 = io_gameIndex == 4'h7 ? cpu_io_dout : _GEN_1175; // @[Main.scala 393:42 MemMap.scala 153:15]
  wire [15:0] eepromMem_din = io_gameIndex == 4'h4 ? cpu_io_dout : _GEN_1368; // @[Main.scala 414:40 MemMap.scala 153:15]
  reg  eeprom_io_serial_cs_r; // @[Reg.scala 35:20]
  wire [23:0] addr_230 = {cpu_io_addr,1'h0}; // @[MemMap.scala 81:25]
  wire  cs_231 = addr_230 >= 24'ha00000 & addr_230 <= 24'ha00000; // @[Util.scala 64:67]
  wire  cs_211 = addr_230 >= 24'hd00000 & addr_230 <= 24'hd00000; // @[Util.scala 64:67]
  wire  cs_179 = addr_230 >= 24'hd00010 & addr_230 <= 24'hd00010; // @[Util.scala 64:67]
  wire  _eepromMem_wr_T_4 = cs_179 & writeStrobe; // @[MemMap.scala 150:20]
  wire  cs_112 = addr_230 >= 24'he00000 & addr_230 <= 24'he00000; // @[Util.scala 64:67]
  wire  cs_26 = addr_230 >= 24'hc00000 & addr_230 <= 24'hc00000; // @[Util.scala 64:67]
  wire  _GEN_236 = io_gameIndex == 4'h0 & (cs_26 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 150:14 MemIO.scala 207:8]
  wire  _GEN_407 = io_gameIndex == 4'h2 ? cs_211 & writeStrobe : _GEN_236; // @[Main.scala 285:42 MemMap.scala 150:14]
  wire  _GEN_572 = io_gameIndex == 4'h1 ? cs_112 & writeStrobe : _GEN_407; // @[Main.scala 306:42 MemMap.scala 150:14]
  wire  _GEN_766 = io_gameIndex == 4'h3 ? cs_112 & writeStrobe : _GEN_572; // @[Main.scala 326:41 MemMap.scala 150:14]
  wire  _GEN_1172 = _cs_T ? cs_179 & writeStrobe : _GEN_766; // @[Main.scala 368:41 MemMap.scala 150:14]
  wire  _GEN_1365 = io_gameIndex == 4'h7 ? cs_211 & writeStrobe : _GEN_1172; // @[Main.scala 393:42 MemMap.scala 150:14]
  wire  eepromMem_wr = io_gameIndex == 4'h4 ? cs_231 & writeStrobe : _GEN_1365; // @[Main.scala 414:40 MemMap.scala 150:14]
  reg  eeprom_io_serial_sck_r; // @[Reg.scala 35:20]
  reg  eeprom_io_serial_sdi_r; // @[Reg.scala 35:20]
  reg  io_gpuMem_layer_0_regs_r_tileSize; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_0_regs_r_enable; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_0_regs_r_flipX; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_0_regs_r_flipY; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_0_regs_r_rowScrollEnable; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_0_regs_r_rowSelectEnable; // @[Reg.scala 19:16]
  reg [8:0] io_gpuMem_layer_0_regs_r_scroll_x; // @[Reg.scala 19:16]
  reg [8:0] io_gpuMem_layer_0_regs_r_scroll_y; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_0_regs_r_1_tileSize; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_0_regs_r_1_enable; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_0_regs_r_1_flipX; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_0_regs_r_1_flipY; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_0_regs_r_1_rowScrollEnable; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_0_regs_r_1_rowSelectEnable; // @[Reg.scala 19:16]
  reg [8:0] io_gpuMem_layer_0_regs_r_1_scroll_x; // @[Reg.scala 19:16]
  reg [8:0] io_gpuMem_layer_0_regs_r_1_scroll_y; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_1_regs_r_tileSize; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_1_regs_r_enable; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_1_regs_r_flipX; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_1_regs_r_flipY; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_1_regs_r_rowScrollEnable; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_1_regs_r_rowSelectEnable; // @[Reg.scala 19:16]
  reg [8:0] io_gpuMem_layer_1_regs_r_scroll_x; // @[Reg.scala 19:16]
  reg [8:0] io_gpuMem_layer_1_regs_r_scroll_y; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_1_regs_r_1_tileSize; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_1_regs_r_1_enable; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_1_regs_r_1_flipX; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_1_regs_r_1_flipY; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_1_regs_r_1_rowScrollEnable; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_1_regs_r_1_rowSelectEnable; // @[Reg.scala 19:16]
  reg [8:0] io_gpuMem_layer_1_regs_r_1_scroll_x; // @[Reg.scala 19:16]
  reg [8:0] io_gpuMem_layer_1_regs_r_1_scroll_y; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_2_regs_r_tileSize; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_2_regs_r_enable; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_2_regs_r_flipX; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_2_regs_r_flipY; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_2_regs_r_rowScrollEnable; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_2_regs_r_rowSelectEnable; // @[Reg.scala 19:16]
  reg [8:0] io_gpuMem_layer_2_regs_r_scroll_x; // @[Reg.scala 19:16]
  reg [8:0] io_gpuMem_layer_2_regs_r_scroll_y; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_2_regs_r_1_tileSize; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_2_regs_r_1_enable; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_2_regs_r_1_flipX; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_2_regs_r_1_flipY; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_2_regs_r_1_rowScrollEnable; // @[Reg.scala 19:16]
  reg  io_gpuMem_layer_2_regs_r_1_rowSelectEnable; // @[Reg.scala 19:16]
  reg [8:0] io_gpuMem_layer_2_regs_r_1_scroll_x; // @[Reg.scala 19:16]
  reg [8:0] io_gpuMem_layer_2_regs_r_1_scroll_y; // @[Reg.scala 19:16]
  reg  REG; // @[Util.scala 165:45]
  wire  _T_1 = ~vBlank & REG; // @[Util.scala 165:35]
  wire  _GEN_60 = _T_1 ? 1'h0 : agalletIrq; // @[Main.scala 213:36 214:16 87:27]
  wire  _GEN_61 = vBlankRising | videoIrq; // @[Main.scala 210:22 211:14 86:25]
  wire  _GEN_62 = vBlankRising | _GEN_60; // @[Main.scala 210:22 212:16]
  reg [21:0] coin1_pulseCounterWrap_value; // @[Counter.scala 40:34]
  wire  coin1_pulseCounterWrap_wrap_wrap = coin1_pulseCounterWrap_value == 22'h30d3ff; // @[Counter.scala 45:24]
  wire [21:0] _coin1_pulseCounterWrap_wrap_value_T_1 = coin1_pulseCounterWrap_value + 22'h1; // @[Counter.scala 46:22]
  reg  coin1_s_enableReg; // @[Util.scala 218:28]
  wire  coin1_pulseCounterWrap = coin1_s_enableReg & coin1_pulseCounterWrap_wrap_wrap; // @[Counter.scala 86:{48,55}]
  reg  coin1_s_REG; // @[Util.scala 158:44]
  wire  _coin1_s_T_1 = io_player_0_coin & ~coin1_s_REG; // @[Util.scala 158:33]
  wire  _GEN_68 = _coin1_s_T_1 | coin1_s_enableReg; // @[Util.scala 218:28 219:{54,66}]
  reg [21:0] coin2_pulseCounterWrap_value; // @[Counter.scala 40:34]
  wire  coin2_pulseCounterWrap_wrap_wrap = coin2_pulseCounterWrap_value == 22'h30d3ff; // @[Counter.scala 45:24]
  wire [21:0] _coin2_pulseCounterWrap_wrap_value_T_1 = coin2_pulseCounterWrap_value + 22'h1; // @[Counter.scala 46:22]
  reg  coin2_s_enableReg; // @[Util.scala 218:28]
  wire  coin2_pulseCounterWrap = coin2_s_enableReg & coin2_pulseCounterWrap_wrap_wrap; // @[Counter.scala 86:{48,55}]
  reg  coin2_s_REG; // @[Util.scala 158:44]
  wire  _coin2_s_T_1 = io_player_1_coin & ~coin2_s_REG; // @[Util.scala 158:33]
  wire  _GEN_75 = _coin2_s_T_1 | coin2_s_enableReg; // @[Util.scala 218:28 219:{54,66}]
  reg [26:0] service_pulseCounterWrap_value; // @[Counter.scala 40:34]
  wire  service_pulseCounterWrap_wrap_wrap = service_pulseCounterWrap_value == 27'h4c4b3ff; // @[Counter.scala 45:24]
  wire [26:0] _service_pulseCounterWrap_wrap_value_T_1 = service_pulseCounterWrap_value + 27'h1; // @[Counter.scala 46:22]
  reg  service_s_enableReg; // @[Util.scala 218:28]
  wire  service_pulseCounterWrap = service_s_enableReg & service_pulseCounterWrap_wrap_wrap; // @[Counter.scala 86:{48,55}]
  reg  service_s_REG; // @[Util.scala 158:44]
  wire  _service_s_T_1 = io_options_service & ~service_s_REG; // @[Util.scala 158:33]
  wire  _GEN_82 = _service_s_T_1 | service_s_enableReg; // @[Util.scala 218:28 219:{54,66}]
  wire  _default1_T = ~service_s_enableReg; // @[Main.scala 447:37]
  wire  _default1_T_1 = ~coin1_s_enableReg; // @[Main.scala 447:47]
  wire  _default1_T_2 = ~io_player_0_start; // @[Main.scala 447:55]
  wire [2:0] _default1_T_4 = ~io_player_0_buttons[2:0]; // @[Main.scala 447:73]
  wire  _default1_T_5 = ~io_player_0_right; // @[Main.scala 447:99]
  wire  _default1_T_6 = ~io_player_0_left; // @[Main.scala 447:117]
  wire  _default1_T_7 = ~io_player_0_down; // @[Main.scala 447:134]
  wire  _default1_T_8 = ~io_player_0_up; // @[Main.scala 447:151]
  wire [15:0] default1 = {6'h3f,_default1_T,_default1_T_1,_default1_T_2,_default1_T_4,_default1_T_5,_default1_T_6,
    _default1_T_7,_default1_T_8}; // @[Cat.scala 33:92]
  wire  _default2_T = ~coin2_s_enableReg; // @[Main.scala 448:66]
  wire  _default2_T_1 = ~io_player_1_start; // @[Main.scala 448:74]
  wire [2:0] _default2_T_3 = ~io_player_1_buttons[2:0]; // @[Main.scala 448:92]
  wire  _default2_T_4 = ~io_player_1_right; // @[Main.scala 448:118]
  wire  _default2_T_5 = ~io_player_1_left; // @[Main.scala 448:136]
  wire  _default2_T_6 = ~io_player_1_down; // @[Main.scala 448:153]
  wire  _default2_T_7 = ~io_player_1_up; // @[Main.scala 448:170]
  wire [15:0] default2 = {4'hf,eeprom_io_serial_sdo,2'h3,_default2_T,_default2_T_1,_default2_T_3,_default2_T_4,
    _default2_T_5,_default2_T_6,_default2_T_7}; // @[Cat.scala 33:92]
  wire [3:0] _left_T_1 = ~io_player_1_buttons; // @[Main.scala 451:26]
  wire [3:0] _left_T_7 = ~io_player_0_buttons; // @[Main.scala 451:119]
  wire [15:0] _left_T_12 = {_left_T_1,_default2_T_4,_default2_T_5,_default2_T_6,_default2_T_7,_left_T_7,_default1_T_5,
    _default1_T_6,_default1_T_7,_default1_T_8}; // @[Cat.scala 33:92]
  wire [7:0] left_lo_1 = {_default1_T_4,_default1_T_5,_default1_T_6,_default1_T_7,_default1_T_8,_default1_T_2}; // @[Cat.scala 33:92]
  wire [15:0] _left_T_27 = {_default2_T_3,_default2_T_4,_default2_T_5,_default2_T_6,_default2_T_7,_default2_T_1,
    left_lo_1}; // @[Cat.scala 33:92]
  wire [15:0] _left_T_29 = 4'h6 == io_gameIndex ? _left_T_12 : default1; // @[Mux.scala 81:58]
  wire [15:0] input0 = 4'h5 == io_gameIndex ? _left_T_27 : _left_T_29; // @[Mux.scala 81:58]
  wire [11:0] _right_T_5 = {6'h3f,_default2_T_1,_default1_T_2,1'h1,_default1_T,_default2_T,_default1_T_1}; // @[Cat.scala 33:92]
  wire [15:0] _right_T_9 = {8'hff,eeprom_io_serial_sdo,4'hf,_default1_T,_default2_T,_default1_T_1}; // @[Cat.scala 33:92]
  wire [15:0] _right_T_11 = 4'h6 == io_gameIndex ? {{4'd0}, _right_T_5} : default2; // @[Mux.scala 81:58]
  wire [15:0] input1 = 4'h5 == io_gameIndex ? _right_T_9 : _right_T_11; // @[Mux.scala 81:58]
  wire  cs_1 = addr_230 >= 24'h110000 & addr_230 <= 24'h1fffff; // @[Util.scala 64:67]
  wire  _GEN_84 = ~cpu_io_as ? 1'h0 : dtackReg; // @[MemMap.scala 226:{19,30} 49:25]
  wire [15:0] _GEN_85 = readStrobe ? 16'h0 : dinReg; // @[MemMap.scala 165:26 166:18 48:23]
  wire [15:0] _GEN_86 = cs_1 ? _GEN_85 : dinReg; // @[MemMap.scala 164:16 48:23]
  wire  _GEN_87 = cs_1 | _GEN_84; // @[MemMap.scala 164:16 170:18]
  wire  cs_2 = addr_230 <= 24'hfffff; // @[Util.scala 64:72]
  wire  _GEN_88 = ~cpu_io_as ? 1'h0 : _GEN_87; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_89 = cs_2 & cpu_io_rw & io_progRom_valid ? io_progRom_dout : _GEN_86; // @[MemMap.scala 130:39 131:16]
  wire  _GEN_90 = cs_2 & cpu_io_rw & io_progRom_valid | _GEN_88; // @[MemMap.scala 130:39 132:18]
  wire  cs_3 = addr_230 >= 24'h100000 & addr_230 <= 24'h10ffff; // @[Util.scala 64:67]
  wire  _GEN_91 = ~cpu_io_as ? 1'h0 : _GEN_90; // @[MemMap.scala 226:{19,30}]
  wire [1:0] _mainRam_io_mask_T = {cpu_io_uds,cpu_io_lds}; // @[MemMap.scala 106:27]
  wire [15:0] _GEN_92 = cs_3 ? mainRam_io_dout : _GEN_89; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_93 = cs_3 | _GEN_91; // @[MemMap.scala 108:16 110:18]
  wire [23:0] offset_3 = addr_230 - 24'h300000; // @[MemMap.scala 84:23]
  wire  cs_4 = addr_230 >= 24'h300000 & addr_230 <= 24'h300003; // @[Util.scala 64:67]
  wire  _GEN_94 = ~cpu_io_as ? 1'h0 : _GEN_93; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_95 = cs_4 ? io_soundCtrl_ymz_dout : _GEN_92; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_96 = cs_4 | _GEN_94; // @[MemMap.scala 108:16 110:18]
  wire  cs_5 = addr_230 >= 24'h400000 & addr_230 <= 24'h40ffff; // @[Util.scala 64:67]
  wire  _GEN_97 = ~cpu_io_as ? 1'h0 : _GEN_96; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_98 = cs_5 ? spriteRam_io_portA_dout : _GEN_95; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_99 = cs_5 | _GEN_97; // @[MemMap.scala 108:16 110:18]
  wire  cs_6 = addr_230 >= 24'h500000 & addr_230 <= 24'h500fff; // @[Util.scala 64:67]
  wire  _GEN_100 = ~cpu_io_as ? 1'h0 : _GEN_99; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_101 = cs_6 ? vram16x16_0_io_portA_dout : _GEN_98; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_102 = cs_6 | _GEN_100; // @[MemMap.scala 108:16 110:18]
  wire  cs_7 = addr_230 >= 24'h501000 & addr_230 <= 24'h5017ff; // @[Util.scala 64:67]
  wire  _GEN_103 = ~cpu_io_as ? 1'h0 : _GEN_102; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_104 = cs_7 ? lineRam_0_io_portA_dout : _GEN_101; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_105 = cs_7 | _GEN_103; // @[MemMap.scala 108:16 110:18]
  wire  cs_8 = addr_230 >= 24'h501800 & addr_230 <= 24'h503fff; // @[Util.scala 64:67]
  wire  _GEN_106 = ~cpu_io_as ? 1'h0 : _GEN_105; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_108 = readStrobe ? tmp : _GEN_104; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_110 = cs_8 ? _GEN_108 : _GEN_104; // @[MemMap.scala 164:16]
  wire  _GEN_112 = cs_8 | _GEN_106; // @[MemMap.scala 164:16 170:18]
  wire  cs_9 = addr_230 >= 24'h504000 & addr_230 <= 24'h507fff; // @[Util.scala 64:67]
  wire  _GEN_113 = ~cpu_io_as ? 1'h0 : _GEN_112; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_114 = cs_9 ? vram8x8_0_io_portA_dout : _GEN_110; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_115 = cs_9 | _GEN_113; // @[MemMap.scala 108:16 110:18]
  wire  cs_10 = addr_230 >= 24'h508000 & addr_230 <= 24'h50ffff; // @[Util.scala 64:67]
  wire  _GEN_116 = ~cpu_io_as ? 1'h0 : _GEN_115; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_1; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_118 = readStrobe ? tmp_1 : _GEN_114; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_120 = cs_10 ? _GEN_118 : _GEN_114; // @[MemMap.scala 164:16]
  wire  _GEN_122 = cs_10 | _GEN_116; // @[MemMap.scala 164:16 170:18]
  wire [23:0] offset_10 = addr_230 - 24'h600000; // @[MemMap.scala 84:23]
  wire  cs_11 = addr_230 >= 24'h600000 & addr_230 <= 24'h600fff; // @[Util.scala 64:67]
  wire  _GEN_123 = ~cpu_io_as ? 1'h0 : _GEN_122; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_124 = cs_11 ? vram16x16_1_io_portA_dout : _GEN_120; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_125 = cs_11 | _GEN_123; // @[MemMap.scala 108:16 110:18]
  wire  cs_12 = addr_230 >= 24'h601000 & addr_230 <= 24'h6017ff; // @[Util.scala 64:67]
  wire  _GEN_126 = ~cpu_io_as ? 1'h0 : _GEN_125; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_127 = cs_12 ? lineRam_1_io_portA_dout : _GEN_124; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_128 = cs_12 | _GEN_126; // @[MemMap.scala 108:16 110:18]
  wire  cs_13 = addr_230 >= 24'h601800 & addr_230 <= 24'h603fff; // @[Util.scala 64:67]
  wire  _GEN_129 = ~cpu_io_as ? 1'h0 : _GEN_128; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_2; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_131 = readStrobe ? tmp_2 : _GEN_127; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_133 = cs_13 ? _GEN_131 : _GEN_127; // @[MemMap.scala 164:16]
  wire  _GEN_135 = cs_13 | _GEN_129; // @[MemMap.scala 164:16 170:18]
  wire  cs_14 = addr_230 >= 24'h604000 & addr_230 <= 24'h607fff; // @[Util.scala 64:67]
  wire  _GEN_136 = ~cpu_io_as ? 1'h0 : _GEN_135; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_137 = cs_14 ? vram8x8_1_io_portA_dout : _GEN_133; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_138 = cs_14 | _GEN_136; // @[MemMap.scala 108:16 110:18]
  wire  cs_15 = addr_230 >= 24'h608000 & addr_230 <= 24'h60ffff; // @[Util.scala 64:67]
  wire  _GEN_139 = ~cpu_io_as ? 1'h0 : _GEN_138; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_3; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_141 = readStrobe ? tmp_3 : _GEN_137; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_143 = cs_15 ? _GEN_141 : _GEN_137; // @[MemMap.scala 164:16]
  wire  _GEN_145 = cs_15 | _GEN_139; // @[MemMap.scala 164:16 170:18]
  wire  cs_16 = addr_230 >= 24'h708000 & addr_230 <= 24'h708fff; // @[Util.scala 64:67]
  wire  _GEN_146 = ~cpu_io_as ? 1'h0 : _GEN_145; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_147 = cs_16 ? paletteRam_io_portA_dout : _GEN_143; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_148 = cs_16 | _GEN_146; // @[MemMap.scala 108:16 110:18]
  wire  cs_17 = addr_230 >= 24'h710c12 & addr_230 <= 24'h710c1f; // @[Util.scala 64:67]
  wire  _GEN_149 = ~cpu_io_as ? 1'h0 : _GEN_148; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_150 = readStrobe ? 16'h0 : _GEN_147; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_151 = cs_17 ? _GEN_150 : _GEN_147; // @[MemMap.scala 164:16]
  wire  _GEN_152 = cs_17 | _GEN_149; // @[MemMap.scala 164:16 170:18]
  wire [23:0] offset_17 = addr_230 - 24'h800000; // @[MemMap.scala 84:23]
  wire  cs_18 = addr_230 >= 24'h800000 & addr_230 <= 24'h800007; // @[Util.scala 64:67]
  wire  _GEN_153 = ~cpu_io_as ? 1'h0 : _GEN_152; // @[MemMap.scala 226:{19,30}]
  wire  dinReg_a = offset_17 == 24'h0 & agalletIrq; // @[Main.scala 219:28]
  wire  _GEN_154 = offset_17 == 24'h4 ? 1'h0 : _GEN_61; // @[Main.scala 222:{26,37}]
  wire  _dinReg_T_2 = ~dinReg_a; // @[Main.scala 224:9]
  wire  _dinReg_T_4 = ~videoIrq; // @[Main.scala 224:17]
  wire [2:0] _dinReg_T_5 = {_dinReg_T_2,1'h1,_dinReg_T_4}; // @[Cat.scala 33:92]
  wire  _GEN_156 = cs_18 & readStrobe ? _GEN_154 : _GEN_61; // @[MemMap.scala 180:30]
  wire [15:0] _GEN_158 = cs_18 & readStrobe ? {{13'd0}, _dinReg_T_5} : _GEN_151; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_159 = cs_18 & readStrobe | _GEN_153; // @[MemMap.scala 180:30 182:18]
  wire  cs_19 = addr_230 >= 24'h800000 & addr_230 <= 24'h80000f; // @[Util.scala 64:67]
  wire  _GEN_160 = ~cpu_io_as ? 1'h0 : _GEN_159; // @[MemMap.scala 226:{19,30}]
  wire  mem_wr = cs_19 & writeStrobe; // @[MemMap.scala 150:20]
  wire  _GEN_161 = cs_19 & _upperWriteStrobe_T_3 | _GEN_160; // @[MemMap.scala 154:{27,38}]
  wire  cs_20 = addr_230 >= 24'h800008 & addr_230 <= 24'h800008; // @[Util.scala 64:67]
  wire  _GEN_162 = ~cpu_io_as ? 1'h0 : _GEN_161; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_163 = cs_20 & writeStrobe | vBlankRising & (_T_260 | pauseReg); // @[MemMap.scala 192:31 Main.scala 232:28 258:68]
  wire  _GEN_164 = cs_20 & writeStrobe | _GEN_162; // @[MemMap.scala 192:31 194:18]
  wire  cs_21 = addr_230 >= 24'h80000a & addr_230 <= 24'h80007f; // @[Util.scala 64:67]
  wire  _GEN_165 = ~cpu_io_as ? 1'h0 : _GEN_164; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_166 = readStrobe ? 16'h0 : _GEN_158; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_167 = cs_21 ? _GEN_166 : _GEN_158; // @[MemMap.scala 164:16]
  wire  _GEN_168 = cs_21 | _GEN_165; // @[MemMap.scala 164:16 170:18]
  wire [23:0] offset_21 = addr_230 - 24'h900000; // @[MemMap.scala 84:23]
  wire  cs_22 = addr_230 >= 24'h900000 & addr_230 <= 24'h900005; // @[Util.scala 64:67]
  wire  _GEN_169 = ~cpu_io_as ? 1'h0 : _GEN_168; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_170 = cs_22 ? layerRegs_0_io_mem_dout : _GEN_167; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_171 = cs_22 | _GEN_169; // @[MemMap.scala 108:16 110:18]
  wire  cs_23 = addr_230 >= 24'ha00000 & addr_230 <= 24'ha00005; // @[Util.scala 64:67]
  wire  _GEN_172 = ~cpu_io_as ? 1'h0 : _GEN_171; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_173 = cs_23 ? layerRegs_1_io_mem_dout : _GEN_170; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_174 = cs_23 | _GEN_172; // @[MemMap.scala 108:16 110:18]
  wire  cs_24 = addr_230 >= 24'hb00000 & addr_230 <= 24'hb00000; // @[Util.scala 64:67]
  wire  _GEN_175 = ~cpu_io_as ? 1'h0 : _GEN_174; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_176 = cs_24 & readStrobe ? input0 : _GEN_173; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_177 = cs_24 & readStrobe | _GEN_175; // @[MemMap.scala 180:30 182:18]
  wire  cs_25 = addr_230 >= 24'hb00002 & addr_230 <= 24'hb00002; // @[Util.scala 64:67]
  wire  _GEN_178 = ~cpu_io_as ? 1'h0 : _GEN_177; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_179 = cs_25 & readStrobe ? input1 : _GEN_176; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_180 = cs_25 & readStrobe | _GEN_178; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_181 = ~cpu_io_as ? 1'h0 : _GEN_180; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_182 = cs_26 & _upperWriteStrobe_T_3 | _GEN_181; // @[MemMap.scala 154:{27,38}]
  wire  _GEN_183 = io_gameIndex == 4'h0 ? _GEN_182 : _GEN_87; // @[Main.scala 267:42]
  wire  _GEN_186 = io_gameIndex == 4'h0 & (cs_2 & readStrobe); // @[Main.scala 267:42 MemMap.scala 128:14 MemIO.scala 83:8]
  wire [15:0] _GEN_188 = io_gameIndex == 4'h0 ? _GEN_179 : _GEN_86; // @[Main.scala 267:42]
  wire  _GEN_189 = io_gameIndex == 4'h0 & (cs_3 & readStrobe); // @[Main.scala 267:42 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_190 = io_gameIndex == 4'h0 & (cs_3 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire [22:0] _GEN_191 = cpu_io_addr; // @[Main.scala 267:42 MemMap.scala 105:16]
  wire  _GEN_194 = io_gameIndex == 4'h0 & (cs_4 & readStrobe); // @[Main.scala 267:42 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_195 = io_gameIndex == 4'h0 & (cs_4 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_197 = io_gameIndex == 4'h0 & (cs_5 & readStrobe); // @[Main.scala 267:42 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_198 = io_gameIndex == 4'h0 & (cs_5 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_200 = io_gameIndex == 4'h0 & (cs_6 & readStrobe); // @[Main.scala 267:42 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_201 = io_gameIndex == 4'h0 & (cs_6 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_203 = io_gameIndex == 4'h0 & (cs_7 & readStrobe); // @[Main.scala 267:42 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_204 = io_gameIndex == 4'h0 & (cs_7 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_206 = io_gameIndex == 4'h0 & (cs_9 & readStrobe); // @[Main.scala 267:42 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_207 = io_gameIndex == 4'h0 & (cs_9 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_209 = io_gameIndex == 4'h0 & (cs_11 & readStrobe); // @[Main.scala 267:42 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_210 = io_gameIndex == 4'h0 & (cs_11 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_212 = io_gameIndex == 4'h0 & (cs_12 & readStrobe); // @[Main.scala 267:42 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_213 = io_gameIndex == 4'h0 & (cs_12 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_215 = io_gameIndex == 4'h0 & (cs_14 & readStrobe); // @[Main.scala 267:42 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_216 = io_gameIndex == 4'h0 & (cs_14 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_218 = io_gameIndex == 4'h0 & (cs_16 & readStrobe); // @[Main.scala 267:42 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_219 = io_gameIndex == 4'h0 & (cs_16 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_222 = io_gameIndex == 4'h0 ? _GEN_156 : _GEN_61; // @[Main.scala 267:42]
  wire  _GEN_225 = io_gameIndex == 4'h0 & mem_wr; // @[Main.scala 267:42 MemIO.scala 305:8 318:8]
  wire [2:0] mem_addr = cpu_io_addr[2:0]; // @[MemIO.scala 303:19 MemMap.scala 151:16]
  wire  _GEN_229 = io_gameIndex == 4'h0 ? _GEN_163 : vBlankRising & (_T_260 | pauseReg); // @[Main.scala 232:28 267:42]
  wire  _GEN_231 = io_gameIndex == 4'h0 & (cs_22 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_234 = io_gameIndex == 4'h0 & (cs_23 & writeStrobe); // @[Main.scala 267:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  cs_27 = addr_230 <= 24'h7ffff; // @[Util.scala 64:72]
  wire  _GEN_238 = ~cpu_io_as ? 1'h0 : _GEN_183; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_239 = cs_27 & cpu_io_rw & io_progRom_valid ? io_progRom_dout : _GEN_188; // @[MemMap.scala 130:39 131:16]
  wire  _GEN_240 = cs_27 & cpu_io_rw & io_progRom_valid | _GEN_238; // @[MemMap.scala 130:39 132:18]
  wire  _GEN_241 = ~cpu_io_as ? 1'h0 : _GEN_240; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_242 = cs_3 ? mainRam_io_dout : _GEN_239; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_243 = cs_3 | _GEN_241; // @[MemMap.scala 108:16 110:18]
  wire  cs_29 = addr_230 >= 24'h200000 & addr_230 <= 24'h200fff; // @[Util.scala 64:67]
  wire  _GEN_244 = ~cpu_io_as ? 1'h0 : _GEN_243; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_245 = cs_29 ? vram16x16_1_io_portA_dout : _GEN_242; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_246 = cs_29 | _GEN_244; // @[MemMap.scala 108:16 110:18]
  wire  cs_30 = addr_230 >= 24'h201000 & addr_230 <= 24'h2017ff; // @[Util.scala 64:67]
  wire  _GEN_247 = ~cpu_io_as ? 1'h0 : _GEN_246; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_248 = cs_30 ? lineRam_1_io_portA_dout : _GEN_245; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_249 = cs_30 | _GEN_247; // @[MemMap.scala 108:16 110:18]
  wire  cs_31 = addr_230 >= 24'h201800 & addr_230 <= 24'h203fff; // @[Util.scala 64:67]
  wire  _GEN_250 = ~cpu_io_as ? 1'h0 : _GEN_249; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_4; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_252 = readStrobe ? tmp_4 : _GEN_248; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_254 = cs_31 ? _GEN_252 : _GEN_248; // @[MemMap.scala 164:16]
  wire  _GEN_256 = cs_31 | _GEN_250; // @[MemMap.scala 164:16 170:18]
  wire  cs_32 = addr_230 >= 24'h204000 & addr_230 <= 24'h207fff; // @[Util.scala 64:67]
  wire  _GEN_257 = ~cpu_io_as ? 1'h0 : _GEN_256; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_258 = cs_32 ? vram8x8_1_io_portA_dout : _GEN_254; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_259 = cs_32 | _GEN_257; // @[MemMap.scala 108:16 110:18]
  wire  cs_33 = addr_230 >= 24'h208000 & addr_230 <= 24'h20ffff; // @[Util.scala 64:67]
  wire  _GEN_260 = ~cpu_io_as ? 1'h0 : _GEN_259; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_5; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_262 = readStrobe ? tmp_5 : _GEN_258; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_264 = cs_33 ? _GEN_262 : _GEN_258; // @[MemMap.scala 164:16]
  wire  _GEN_266 = cs_33 | _GEN_260; // @[MemMap.scala 164:16 170:18]
  wire  cs_34 = addr_230 >= 24'h300000 & addr_230 <= 24'h300fff; // @[Util.scala 64:67]
  wire  _GEN_267 = ~cpu_io_as ? 1'h0 : _GEN_266; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_268 = cs_34 ? vram16x16_0_io_portA_dout : _GEN_264; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_269 = cs_34 | _GEN_267; // @[MemMap.scala 108:16 110:18]
  wire  cs_35 = addr_230 >= 24'h301000 & addr_230 <= 24'h3017ff; // @[Util.scala 64:67]
  wire  _GEN_270 = ~cpu_io_as ? 1'h0 : _GEN_269; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_271 = cs_35 ? lineRam_0_io_portA_dout : _GEN_268; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_272 = cs_35 | _GEN_270; // @[MemMap.scala 108:16 110:18]
  wire  cs_36 = addr_230 >= 24'h301800 & addr_230 <= 24'h303fff; // @[Util.scala 64:67]
  wire  _GEN_273 = ~cpu_io_as ? 1'h0 : _GEN_272; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_6; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_275 = readStrobe ? tmp_6 : _GEN_271; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_277 = cs_36 ? _GEN_275 : _GEN_271; // @[MemMap.scala 164:16]
  wire  _GEN_279 = cs_36 | _GEN_273; // @[MemMap.scala 164:16 170:18]
  wire  cs_37 = addr_230 >= 24'h304000 & addr_230 <= 24'h307fff; // @[Util.scala 64:67]
  wire  _GEN_280 = ~cpu_io_as ? 1'h0 : _GEN_279; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_281 = cs_37 ? vram8x8_0_io_portA_dout : _GEN_277; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_282 = cs_37 | _GEN_280; // @[MemMap.scala 108:16 110:18]
  wire  cs_38 = addr_230 >= 24'h308000 & addr_230 <= 24'h30ffff; // @[Util.scala 64:67]
  wire  _GEN_283 = ~cpu_io_as ? 1'h0 : _GEN_282; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_7; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_285 = readStrobe ? tmp_7 : _GEN_281; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_287 = cs_38 ? _GEN_285 : _GEN_281; // @[MemMap.scala 164:16]
  wire  _GEN_289 = cs_38 | _GEN_283; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_290 = ~cpu_io_as ? 1'h0 : _GEN_289; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_291 = cs_5 ? vram8x8_2_io_portA_dout : _GEN_287; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_292 = cs_5 | _GEN_290; // @[MemMap.scala 108:16 110:18]
  wire  cs_40 = addr_230 >= 24'h500000 & addr_230 <= 24'h50ffff; // @[Util.scala 64:67]
  wire  _GEN_293 = ~cpu_io_as ? 1'h0 : _GEN_292; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_294 = cs_40 ? spriteRam_io_portA_dout : _GEN_291; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_295 = cs_40 | _GEN_293; // @[MemMap.scala 108:16 110:18]
  wire  cs_41 = addr_230 >= 24'h600000 & addr_230 <= 24'h600005; // @[Util.scala 64:67]
  wire  _GEN_296 = ~cpu_io_as ? 1'h0 : _GEN_295; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_297 = cs_41 ? layerRegs_1_io_mem_dout : _GEN_294; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_298 = cs_41 | _GEN_296; // @[MemMap.scala 108:16 110:18]
  wire  cs_42 = addr_230 >= 24'h700000 & addr_230 <= 24'h700005; // @[Util.scala 64:67]
  wire  _GEN_299 = ~cpu_io_as ? 1'h0 : _GEN_298; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_300 = cs_42 ? layerRegs_0_io_mem_dout : _GEN_297; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_301 = cs_42 | _GEN_299; // @[MemMap.scala 108:16 110:18]
  wire  cs_43 = addr_230 >= 24'h800000 & addr_230 <= 24'h800005; // @[Util.scala 64:67]
  wire  _GEN_302 = ~cpu_io_as ? 1'h0 : _GEN_301; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_303 = cs_43 ? layerRegs_2_io_mem_dout : _GEN_300; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_304 = cs_43 | _GEN_302; // @[MemMap.scala 108:16 110:18]
  wire  cs_44 = addr_230 >= 24'h900000 & addr_230 <= 24'h900007; // @[Util.scala 64:67]
  wire  _GEN_305 = ~cpu_io_as ? 1'h0 : _GEN_304; // @[MemMap.scala 226:{19,30}]
  wire  dinReg_a_1 = offset_21 == 24'h0 & agalletIrq; // @[Main.scala 219:28]
  wire  _GEN_306 = offset_21 == 24'h4 ? 1'h0 : _GEN_222; // @[Main.scala 222:{26,37}]
  wire  _dinReg_T_8 = ~dinReg_a_1; // @[Main.scala 224:9]
  wire [2:0] _dinReg_T_11 = {_dinReg_T_8,1'h1,_dinReg_T_4}; // @[Cat.scala 33:92]
  wire  _GEN_308 = cs_44 & readStrobe ? _GEN_306 : _GEN_222; // @[MemMap.scala 180:30]
  wire [15:0] _GEN_310 = cs_44 & readStrobe ? {{13'd0}, _dinReg_T_11} : _GEN_303; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_311 = cs_44 & readStrobe | _GEN_305; // @[MemMap.scala 180:30 182:18]
  wire  cs_45 = addr_230 >= 24'h900000 & addr_230 <= 24'h90000f; // @[Util.scala 64:67]
  wire  _GEN_312 = ~cpu_io_as ? 1'h0 : _GEN_311; // @[MemMap.scala 226:{19,30}]
  wire  mem_1_wr = cs_45 & writeStrobe; // @[MemMap.scala 150:20]
  wire  _GEN_313 = cs_45 & _upperWriteStrobe_T_3 | _GEN_312; // @[MemMap.scala 154:{27,38}]
  wire  cs_46 = addr_230 >= 24'h900008 & addr_230 <= 24'h900008; // @[Util.scala 64:67]
  wire  _GEN_314 = ~cpu_io_as ? 1'h0 : _GEN_313; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_315 = cs_46 & writeStrobe | _GEN_229; // @[MemMap.scala 192:31 Main.scala 258:68]
  wire  _GEN_316 = cs_46 & writeStrobe | _GEN_314; // @[MemMap.scala 192:31 194:18]
  wire  cs_47 = addr_230 >= 24'h90000a & addr_230 <= 24'h90007f; // @[Util.scala 64:67]
  wire  _GEN_317 = ~cpu_io_as ? 1'h0 : _GEN_316; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_318 = readStrobe ? 16'h0 : _GEN_310; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_319 = cs_47 ? _GEN_318 : _GEN_310; // @[MemMap.scala 164:16]
  wire  _GEN_320 = cs_47 | _GEN_317; // @[MemMap.scala 164:16 170:18]
  wire  cs_48 = addr_230 >= 24'ha08000 & addr_230 <= 24'ha08fff; // @[Util.scala 64:67]
  wire  _GEN_321 = ~cpu_io_as ? 1'h0 : _GEN_320; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_322 = cs_48 ? paletteRam_io_portA_dout : _GEN_319; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_323 = cs_48 | _GEN_321; // @[MemMap.scala 108:16 110:18]
  wire  cs_49 = addr_230 >= 24'hb00000 & addr_230 <= 24'hb00003; // @[Util.scala 64:67]
  wire  _GEN_324 = ~cpu_io_as ? 1'h0 : _GEN_323; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_325 = cs_49 ? io_soundCtrl_oki_0_dout : _GEN_322; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_326 = cs_49 | _GEN_324; // @[MemMap.scala 108:16 110:18]
  wire  cs_50 = addr_230 >= 24'hb00010 & addr_230 <= 24'hb00013; // @[Util.scala 64:67]
  wire  _GEN_327 = ~cpu_io_as ? 1'h0 : _GEN_326; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_328 = cs_50 ? io_soundCtrl_oki_1_dout : _GEN_325; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_329 = cs_50 | _GEN_327; // @[MemMap.scala 108:16 110:18]
  wire  cs_51 = addr_230 >= 24'hb00020 & addr_230 <= 24'hb0002f; // @[Util.scala 64:67]
  wire  _GEN_330 = ~cpu_io_as ? 1'h0 : _GEN_329; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_331 = cs_51 & _upperWriteStrobe_T_3 | _GEN_330; // @[MemMap.scala 154:{27,38}]
  wire  _GEN_332 = ~cpu_io_as ? 1'h0 : _GEN_331; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_333 = cs_26 & readStrobe ? input0 : _GEN_328; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_334 = cs_26 & readStrobe | _GEN_332; // @[MemMap.scala 180:30 182:18]
  wire  cs_53 = addr_230 >= 24'hc00002 & addr_230 <= 24'hc00002; // @[Util.scala 64:67]
  wire  _GEN_335 = ~cpu_io_as ? 1'h0 : _GEN_334; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_336 = cs_53 & readStrobe ? input1 : _GEN_333; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_337 = cs_53 & readStrobe | _GEN_335; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_338 = ~cpu_io_as ? 1'h0 : _GEN_337; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_339 = cs_211 & _upperWriteStrobe_T_3 | _GEN_338; // @[MemMap.scala 154:{27,38}]
  wire  _GEN_340 = io_gameIndex == 4'h2 ? _GEN_339 : _GEN_183; // @[Main.scala 285:42]
  wire  _GEN_343 = io_gameIndex == 4'h2 ? cs_27 & readStrobe : _GEN_186; // @[Main.scala 285:42 MemMap.scala 128:14]
  wire [23:0] _GEN_344 = io_gameIndex == 4'h2 ? addr_230 : addr_230; // @[Main.scala 285:42 MemMap.scala 129:16]
  wire [15:0] _GEN_345 = io_gameIndex == 4'h2 ? _GEN_336 : _GEN_188; // @[Main.scala 285:42]
  wire  _GEN_346 = io_gameIndex == 4'h2 ? cs_3 & readStrobe : _GEN_189; // @[Main.scala 285:42 MemMap.scala 103:14]
  wire  _GEN_347 = io_gameIndex == 4'h2 ? cs_3 & writeStrobe : _GEN_190; // @[Main.scala 285:42 MemMap.scala 104:14]
  wire [22:0] _GEN_348 = io_gameIndex == 4'h2 ? cpu_io_addr : _GEN_191; // @[Main.scala 285:42 MemMap.scala 105:16]
  wire [1:0] _GEN_349 = io_gameIndex == 4'h2 ? _mainRam_io_mask_T : _mainRam_io_mask_T; // @[Main.scala 285:42 MemMap.scala 106:16]
  wire  _GEN_351 = io_gameIndex == 4'h2 ? cs_29 & readStrobe : _GEN_209; // @[Main.scala 285:42 MemMap.scala 103:14]
  wire  _GEN_352 = io_gameIndex == 4'h2 ? cs_29 & writeStrobe : _GEN_210; // @[Main.scala 285:42 MemMap.scala 104:14]
  wire  _GEN_354 = io_gameIndex == 4'h2 ? cs_30 & readStrobe : _GEN_212; // @[Main.scala 285:42 MemMap.scala 103:14]
  wire  _GEN_355 = io_gameIndex == 4'h2 ? cs_30 & writeStrobe : _GEN_213; // @[Main.scala 285:42 MemMap.scala 104:14]
  wire  _GEN_357 = io_gameIndex == 4'h2 ? cs_32 & readStrobe : _GEN_215; // @[Main.scala 285:42 MemMap.scala 103:14]
  wire  _GEN_358 = io_gameIndex == 4'h2 ? cs_32 & writeStrobe : _GEN_216; // @[Main.scala 285:42 MemMap.scala 104:14]
  wire  _GEN_360 = io_gameIndex == 4'h2 ? cs_34 & readStrobe : _GEN_200; // @[Main.scala 285:42 MemMap.scala 103:14]
  wire  _GEN_361 = io_gameIndex == 4'h2 ? cs_34 & writeStrobe : _GEN_201; // @[Main.scala 285:42 MemMap.scala 104:14]
  wire  _GEN_363 = io_gameIndex == 4'h2 ? cs_35 & readStrobe : _GEN_203; // @[Main.scala 285:42 MemMap.scala 103:14]
  wire  _GEN_364 = io_gameIndex == 4'h2 ? cs_35 & writeStrobe : _GEN_204; // @[Main.scala 285:42 MemMap.scala 104:14]
  wire  _GEN_366 = io_gameIndex == 4'h2 ? cs_37 & readStrobe : _GEN_206; // @[Main.scala 285:42 MemMap.scala 103:14]
  wire  _GEN_367 = io_gameIndex == 4'h2 ? cs_37 & writeStrobe : _GEN_207; // @[Main.scala 285:42 MemMap.scala 104:14]
  wire  _GEN_369 = io_gameIndex == 4'h2 & (cs_5 & readStrobe); // @[Main.scala 285:42 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_370 = io_gameIndex == 4'h2 & (cs_5 & writeStrobe); // @[Main.scala 285:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_374 = io_gameIndex == 4'h2 ? cs_40 & readStrobe : _GEN_197; // @[Main.scala 285:42 MemMap.scala 103:14]
  wire  _GEN_375 = io_gameIndex == 4'h2 ? cs_40 & writeStrobe : _GEN_198; // @[Main.scala 285:42 MemMap.scala 104:14]
  wire  _GEN_378 = io_gameIndex == 4'h2 ? cs_41 & writeStrobe : _GEN_234; // @[Main.scala 285:42 MemMap.scala 104:14]
  wire  _GEN_381 = io_gameIndex == 4'h2 ? cs_42 & writeStrobe : _GEN_231; // @[Main.scala 285:42 MemMap.scala 104:14]
  wire  _GEN_384 = io_gameIndex == 4'h2 & (cs_43 & writeStrobe); // @[Main.scala 285:42 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_387 = io_gameIndex == 4'h2 ? _GEN_308 : _GEN_222; // @[Main.scala 285:42]
  wire  _GEN_390 = io_gameIndex == 4'h2 ? mem_1_wr : _GEN_225; // @[Main.scala 285:42 MemIO.scala 305:8]
  wire [2:0] _GEN_391 = io_gameIndex == 4'h2 ? mem_addr : mem_addr; // @[Main.scala 285:42 MemIO.scala 306:10]
  wire [15:0] _GEN_393 = io_gameIndex == 4'h2 ? _GEN_193 : _GEN_193; // @[Main.scala 285:42 MemIO.scala 308:9]
  wire  _GEN_394 = io_gameIndex == 4'h2 ? _GEN_315 : _GEN_229; // @[Main.scala 285:42]
  wire  _GEN_395 = io_gameIndex == 4'h2 ? cs_48 & readStrobe : _GEN_218; // @[Main.scala 285:42 MemMap.scala 103:14]
  wire  _GEN_396 = io_gameIndex == 4'h2 ? cs_48 & writeStrobe : _GEN_219; // @[Main.scala 285:42 MemMap.scala 104:14]
  wire [10:0] _GEN_397 = io_gameIndex == 4'h2 ? cpu_io_addr[10:0] : cpu_io_addr[10:0]; // @[Main.scala 285:42 MemMap.scala 105:16]
  wire  _GEN_409 = ~cpu_io_as ? 1'h0 : _GEN_340; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_410 = cs_2 & cpu_io_rw & io_progRom_valid ? io_progRom_dout : _GEN_345; // @[MemMap.scala 130:39 131:16]
  wire  _GEN_411 = cs_2 & cpu_io_rw & io_progRom_valid | _GEN_409; // @[MemMap.scala 130:39 132:18]
  wire  _GEN_412 = ~cpu_io_as ? 1'h0 : _GEN_411; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_413 = cs_3 ? mainRam_io_dout : _GEN_410; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_414 = cs_3 | _GEN_412; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_415 = ~cpu_io_as ? 1'h0 : _GEN_414; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_416 = cs_4 ? io_soundCtrl_ymz_dout : _GEN_413; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_417 = cs_4 | _GEN_415; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_418 = ~cpu_io_as ? 1'h0 : _GEN_417; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_419 = cs_5 ? spriteRam_io_portA_dout : _GEN_416; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_420 = cs_5 | _GEN_418; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_421 = ~cpu_io_as ? 1'h0 : _GEN_420; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_422 = cs_6 ? vram16x16_0_io_portA_dout : _GEN_419; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_423 = cs_6 | _GEN_421; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_424 = ~cpu_io_as ? 1'h0 : _GEN_423; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_425 = cs_7 ? lineRam_0_io_portA_dout : _GEN_422; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_426 = cs_7 | _GEN_424; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_427 = ~cpu_io_as ? 1'h0 : _GEN_426; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_8; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_429 = readStrobe ? tmp_8 : _GEN_425; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_431 = cs_8 ? _GEN_429 : _GEN_425; // @[MemMap.scala 164:16]
  wire  _GEN_433 = cs_8 | _GEN_427; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_434 = ~cpu_io_as ? 1'h0 : _GEN_433; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_435 = cs_9 ? vram8x8_0_io_portA_dout : _GEN_431; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_436 = cs_9 | _GEN_434; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_437 = ~cpu_io_as ? 1'h0 : _GEN_436; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_9; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_439 = readStrobe ? tmp_9 : _GEN_435; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_441 = cs_10 ? _GEN_439 : _GEN_435; // @[MemMap.scala 164:16]
  wire  _GEN_443 = cs_10 | _GEN_437; // @[MemMap.scala 164:16 170:18]
  wire  cs_64 = addr_230 >= 24'h5fff00 & addr_230 <= 24'h5fffff; // @[Util.scala 64:67]
  wire  _GEN_444 = ~cpu_io_as ? 1'h0 : _GEN_443; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_445 = cs_64 & writeStrobe | _GEN_444; // @[MemMap.scala 192:31 194:18]
  wire  _GEN_446 = ~cpu_io_as ? 1'h0 : _GEN_445; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_447 = cs_11 ? vram16x16_1_io_portA_dout : _GEN_441; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_448 = cs_11 | _GEN_446; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_449 = ~cpu_io_as ? 1'h0 : _GEN_448; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_450 = cs_12 ? lineRam_1_io_portA_dout : _GEN_447; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_451 = cs_12 | _GEN_449; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_452 = ~cpu_io_as ? 1'h0 : _GEN_451; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_10; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_454 = readStrobe ? tmp_10 : _GEN_450; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_456 = cs_13 ? _GEN_454 : _GEN_450; // @[MemMap.scala 164:16]
  wire  _GEN_458 = cs_13 | _GEN_452; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_459 = ~cpu_io_as ? 1'h0 : _GEN_458; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_460 = cs_14 ? vram8x8_1_io_portA_dout : _GEN_456; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_461 = cs_14 | _GEN_459; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_462 = ~cpu_io_as ? 1'h0 : _GEN_461; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_11; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_464 = readStrobe ? tmp_11 : _GEN_460; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_466 = cs_15 ? _GEN_464 : _GEN_460; // @[MemMap.scala 164:16]
  wire  _GEN_468 = cs_15 | _GEN_462; // @[MemMap.scala 164:16 170:18]
  wire  cs_70 = addr_230 >= 24'h700000 & addr_230 <= 24'h70ffff; // @[Util.scala 64:67]
  wire  _GEN_469 = ~cpu_io_as ? 1'h0 : _GEN_468; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_470 = cs_70 ? vram8x8_2_io_portA_dout : _GEN_466; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_471 = cs_70 | _GEN_469; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_472 = ~cpu_io_as ? 1'h0 : _GEN_471; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_473 = offset_17 == 24'h4 ? 1'h0 : _GEN_387; // @[Main.scala 222:{26,37}]
  wire  _GEN_475 = cs_18 & readStrobe ? _GEN_473 : _GEN_387; // @[MemMap.scala 180:30]
  wire [15:0] _GEN_477 = cs_18 & readStrobe ? {{13'd0}, _dinReg_T_5} : _GEN_470; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_478 = cs_18 & readStrobe | _GEN_472; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_479 = ~cpu_io_as ? 1'h0 : _GEN_478; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_480 = cs_19 & _upperWriteStrobe_T_3 | _GEN_479; // @[MemMap.scala 154:{27,38}]
  wire  _GEN_481 = ~cpu_io_as ? 1'h0 : _GEN_480; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_482 = cs_20 & writeStrobe | _GEN_394; // @[MemMap.scala 192:31 Main.scala 258:68]
  wire  _GEN_483 = cs_20 & writeStrobe | _GEN_481; // @[MemMap.scala 192:31 194:18]
  wire  _GEN_484 = ~cpu_io_as ? 1'h0 : _GEN_483; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_485 = readStrobe ? 16'h0 : _GEN_477; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_486 = cs_21 ? _GEN_485 : _GEN_477; // @[MemMap.scala 164:16]
  wire  _GEN_487 = cs_21 | _GEN_484; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_488 = ~cpu_io_as ? 1'h0 : _GEN_487; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_489 = cs_22 ? layerRegs_0_io_mem_dout : _GEN_486; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_490 = cs_22 | _GEN_488; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_491 = ~cpu_io_as ? 1'h0 : _GEN_490; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_492 = cs_23 ? layerRegs_1_io_mem_dout : _GEN_489; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_493 = cs_23 | _GEN_491; // @[MemMap.scala 108:16 110:18]
  wire  cs_77 = addr_230 >= 24'hb00000 & addr_230 <= 24'hb00005; // @[Util.scala 64:67]
  wire  _GEN_494 = ~cpu_io_as ? 1'h0 : _GEN_493; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_495 = cs_77 ? layerRegs_2_io_mem_dout : _GEN_492; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_496 = cs_77 | _GEN_494; // @[MemMap.scala 108:16 110:18]
  wire  cs_78 = addr_230 >= 24'hc00000 & addr_230 <= 24'hc0ffff; // @[Util.scala 64:67]
  wire  _GEN_497 = ~cpu_io_as ? 1'h0 : _GEN_496; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_498 = cs_78 ? paletteRam_io_portA_dout : _GEN_495; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_499 = cs_78 | _GEN_497; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_500 = ~cpu_io_as ? 1'h0 : _GEN_499; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_501 = cs_211 & readStrobe ? input0 : _GEN_498; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_502 = cs_211 & readStrobe | _GEN_500; // @[MemMap.scala 180:30 182:18]
  wire  cs_80 = addr_230 >= 24'hd00002 & addr_230 <= 24'hd00002; // @[Util.scala 64:67]
  wire  _GEN_503 = ~cpu_io_as ? 1'h0 : _GEN_502; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_504 = cs_80 & readStrobe ? input1 : _GEN_501; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_505 = cs_80 & readStrobe | _GEN_503; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_506 = ~cpu_io_as ? 1'h0 : _GEN_505; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_507 = cs_112 & _upperWriteStrobe_T_3 | _GEN_506; // @[MemMap.scala 154:{27,38}]
  wire  _GEN_508 = io_gameIndex == 4'h1 ? _GEN_507 : _GEN_340; // @[Main.scala 306:42]
  wire  _GEN_511 = io_gameIndex == 4'h1 ? cs_2 & readStrobe : _GEN_343; // @[Main.scala 306:42 MemMap.scala 128:14]
  wire [23:0] _GEN_512 = io_gameIndex == 4'h1 ? addr_230 : _GEN_344; // @[Main.scala 306:42 MemMap.scala 129:16]
  wire [15:0] _GEN_513 = io_gameIndex == 4'h1 ? _GEN_504 : _GEN_345; // @[Main.scala 306:42]
  wire  _GEN_514 = io_gameIndex == 4'h1 ? cs_3 & readStrobe : _GEN_346; // @[Main.scala 306:42 MemMap.scala 103:14]
  wire  _GEN_515 = io_gameIndex == 4'h1 ? cs_3 & writeStrobe : _GEN_347; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire [22:0] _GEN_516 = io_gameIndex == 4'h1 ? cpu_io_addr : _GEN_348; // @[Main.scala 306:42 MemMap.scala 105:16]
  wire [1:0] _GEN_517 = io_gameIndex == 4'h1 ? _mainRam_io_mask_T : _GEN_349; // @[Main.scala 306:42 MemMap.scala 106:16]
  wire  _GEN_519 = io_gameIndex == 4'h1 ? cs_4 & readStrobe : _GEN_194; // @[Main.scala 306:42 MemMap.scala 103:14]
  wire  _GEN_520 = io_gameIndex == 4'h1 ? cs_4 & writeStrobe : _GEN_195; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire [22:0] _GEN_521 = io_gameIndex == 4'h1 ? cpu_io_addr : _GEN_191; // @[Main.scala 306:42 MemMap.scala 105:16]
  wire [1:0] _GEN_522 = io_gameIndex == 4'h1 ? _mainRam_io_mask_T : _mainRam_io_mask_T; // @[Main.scala 306:42 MemMap.scala 106:16]
  wire [15:0] _GEN_523 = io_gameIndex == 4'h1 ? cpu_io_dout : _GEN_193; // @[Main.scala 306:42 MemMap.scala 107:15]
  wire  _GEN_524 = io_gameIndex == 4'h1 ? cs_5 & readStrobe : _GEN_374; // @[Main.scala 306:42 MemMap.scala 103:14]
  wire  _GEN_525 = io_gameIndex == 4'h1 ? cs_5 & writeStrobe : _GEN_375; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire  _GEN_527 = io_gameIndex == 4'h1 ? cs_6 & readStrobe : _GEN_360; // @[Main.scala 306:42 MemMap.scala 103:14]
  wire  _GEN_528 = io_gameIndex == 4'h1 ? cs_6 & writeStrobe : _GEN_361; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire  _GEN_530 = io_gameIndex == 4'h1 ? cs_7 & readStrobe : _GEN_363; // @[Main.scala 306:42 MemMap.scala 103:14]
  wire  _GEN_531 = io_gameIndex == 4'h1 ? cs_7 & writeStrobe : _GEN_364; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire  _GEN_533 = io_gameIndex == 4'h1 ? cs_9 & readStrobe : _GEN_366; // @[Main.scala 306:42 MemMap.scala 103:14]
  wire  _GEN_534 = io_gameIndex == 4'h1 ? cs_9 & writeStrobe : _GEN_367; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire  _GEN_536 = io_gameIndex == 4'h1 ? cs_11 & readStrobe : _GEN_351; // @[Main.scala 306:42 MemMap.scala 103:14]
  wire  _GEN_537 = io_gameIndex == 4'h1 ? cs_11 & writeStrobe : _GEN_352; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire  _GEN_539 = io_gameIndex == 4'h1 ? cs_12 & readStrobe : _GEN_354; // @[Main.scala 306:42 MemMap.scala 103:14]
  wire  _GEN_540 = io_gameIndex == 4'h1 ? cs_12 & writeStrobe : _GEN_355; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire  _GEN_542 = io_gameIndex == 4'h1 ? cs_14 & readStrobe : _GEN_357; // @[Main.scala 306:42 MemMap.scala 103:14]
  wire  _GEN_543 = io_gameIndex == 4'h1 ? cs_14 & writeStrobe : _GEN_358; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire  _GEN_545 = io_gameIndex == 4'h1 ? cs_70 & readStrobe : _GEN_369; // @[Main.scala 306:42 MemMap.scala 103:14]
  wire  _GEN_546 = io_gameIndex == 4'h1 ? cs_70 & writeStrobe : _GEN_370; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire [12:0] _GEN_547 = io_gameIndex == 4'h1 ? cpu_io_addr[12:0] : cpu_io_addr[12:0]; // @[Main.scala 306:42 MemMap.scala 105:16]
  wire  _GEN_550 = io_gameIndex == 4'h1 ? _GEN_475 : _GEN_387; // @[Main.scala 306:42]
  wire  _GEN_553 = io_gameIndex == 4'h1 ? mem_wr : _GEN_390; // @[Main.scala 306:42 MemIO.scala 305:8]
  wire [2:0] _GEN_554 = io_gameIndex == 4'h1 ? mem_addr : _GEN_391; // @[Main.scala 306:42 MemIO.scala 306:10]
  wire [15:0] _GEN_556 = io_gameIndex == 4'h1 ? _GEN_193 : _GEN_393; // @[Main.scala 306:42 MemIO.scala 308:9]
  wire  _GEN_557 = io_gameIndex == 4'h1 ? _GEN_482 : _GEN_394; // @[Main.scala 306:42]
  wire  _GEN_559 = io_gameIndex == 4'h1 ? cs_22 & writeStrobe : _GEN_381; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire  _GEN_562 = io_gameIndex == 4'h1 ? cs_23 & writeStrobe : _GEN_378; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire  _GEN_565 = io_gameIndex == 4'h1 ? cs_77 & writeStrobe : _GEN_384; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire  _GEN_568 = io_gameIndex == 4'h1 ? cs_78 & readStrobe : _GEN_395; // @[Main.scala 306:42 MemMap.scala 103:14]
  wire  _GEN_569 = io_gameIndex == 4'h1 ? cs_78 & writeStrobe : _GEN_396; // @[Main.scala 306:42 MemMap.scala 104:14]
  wire [22:0] _GEN_570 = io_gameIndex == 4'h1 ? cpu_io_addr : {{12'd0}, _GEN_397}; // @[Main.scala 306:42 MemMap.scala 105:16]
  wire  _GEN_574 = ~cpu_io_as ? 1'h0 : _GEN_508; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_575 = cs_2 & cpu_io_rw & io_progRom_valid ? io_progRom_dout : _GEN_513; // @[MemMap.scala 130:39 131:16]
  wire  _GEN_576 = cs_2 & cpu_io_rw & io_progRom_valid | _GEN_574; // @[MemMap.scala 130:39 132:18]
  wire  _GEN_577 = ~cpu_io_as ? 1'h0 : _GEN_576; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_578 = cs_3 ? mainRam_io_dout : _GEN_575; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_579 = cs_3 | _GEN_577; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_580 = ~cpu_io_as ? 1'h0 : _GEN_579; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_581 = cs_4 ? io_soundCtrl_ymz_dout : _GEN_578; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_582 = cs_4 | _GEN_580; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_583 = ~cpu_io_as ? 1'h0 : _GEN_582; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_584 = cs_5 ? spriteRam_io_portA_dout : _GEN_581; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_585 = cs_5 | _GEN_583; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_586 = ~cpu_io_as ? 1'h0 : _GEN_585; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_587 = cs_6 ? vram16x16_0_io_portA_dout : _GEN_584; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_588 = cs_6 | _GEN_586; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_589 = ~cpu_io_as ? 1'h0 : _GEN_588; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_590 = cs_7 ? lineRam_0_io_portA_dout : _GEN_587; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_591 = cs_7 | _GEN_589; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_592 = ~cpu_io_as ? 1'h0 : _GEN_591; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_12; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_594 = readStrobe ? tmp_12 : _GEN_590; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_596 = cs_8 ? _GEN_594 : _GEN_590; // @[MemMap.scala 164:16]
  wire  _GEN_598 = cs_8 | _GEN_592; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_599 = ~cpu_io_as ? 1'h0 : _GEN_598; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_600 = cs_9 ? vram8x8_0_io_portA_dout : _GEN_596; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_601 = cs_9 | _GEN_599; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_602 = ~cpu_io_as ? 1'h0 : _GEN_601; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_13; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_604 = readStrobe ? tmp_13 : _GEN_600; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_606 = cs_10 ? _GEN_604 : _GEN_600; // @[MemMap.scala 164:16]
  wire  _GEN_608 = cs_10 | _GEN_602; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_609 = ~cpu_io_as ? 1'h0 : _GEN_608; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_610 = cs_11 ? vram16x16_1_io_portA_dout : _GEN_606; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_611 = cs_11 | _GEN_609; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_612 = ~cpu_io_as ? 1'h0 : _GEN_611; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_613 = cs_12 ? lineRam_1_io_portA_dout : _GEN_610; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_614 = cs_12 | _GEN_612; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_615 = ~cpu_io_as ? 1'h0 : _GEN_614; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_14; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_617 = readStrobe ? tmp_14 : _GEN_613; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_619 = cs_13 ? _GEN_617 : _GEN_613; // @[MemMap.scala 164:16]
  wire  _GEN_621 = cs_13 | _GEN_615; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_622 = ~cpu_io_as ? 1'h0 : _GEN_621; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_623 = cs_14 ? vram8x8_1_io_portA_dout : _GEN_619; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_624 = cs_14 | _GEN_622; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_625 = ~cpu_io_as ? 1'h0 : _GEN_624; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_15; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_627 = readStrobe ? tmp_15 : _GEN_623; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_629 = cs_15 ? _GEN_627 : _GEN_623; // @[MemMap.scala 164:16]
  wire  _GEN_631 = cs_15 | _GEN_625; // @[MemMap.scala 164:16 170:18]
  wire  cs_96 = addr_230 >= 24'h700000 & addr_230 <= 24'h700fff; // @[Util.scala 64:67]
  wire  _GEN_632 = ~cpu_io_as ? 1'h0 : _GEN_631; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_633 = cs_96 ? vram16x16_2_io_portA_dout : _GEN_629; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_634 = cs_96 | _GEN_632; // @[MemMap.scala 108:16 110:18]
  wire  cs_97 = addr_230 >= 24'h701000 & addr_230 <= 24'h7017ff; // @[Util.scala 64:67]
  wire  _GEN_635 = ~cpu_io_as ? 1'h0 : _GEN_634; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_636 = cs_97 ? lineRam_2_io_portA_dout : _GEN_633; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_637 = cs_97 | _GEN_635; // @[MemMap.scala 108:16 110:18]
  wire  cs_98 = addr_230 >= 24'h701800 & addr_230 <= 24'h703fff; // @[Util.scala 64:67]
  wire  _GEN_638 = ~cpu_io_as ? 1'h0 : _GEN_637; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_16; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_640 = readStrobe ? tmp_16 : _GEN_636; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_642 = cs_98 ? _GEN_640 : _GEN_636; // @[MemMap.scala 164:16]
  wire  _GEN_644 = cs_98 | _GEN_638; // @[MemMap.scala 164:16 170:18]
  wire  cs_99 = addr_230 >= 24'h704000 & addr_230 <= 24'h707fff; // @[Util.scala 64:67]
  wire  _GEN_645 = ~cpu_io_as ? 1'h0 : _GEN_644; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_646 = cs_99 ? vram8x8_2_io_portA_dout : _GEN_642; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_647 = cs_99 | _GEN_645; // @[MemMap.scala 108:16 110:18]
  wire  cs_100 = addr_230 >= 24'h708000 & addr_230 <= 24'h70ffff; // @[Util.scala 64:67]
  wire  _GEN_648 = ~cpu_io_as ? 1'h0 : _GEN_647; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_17; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_650 = readStrobe ? tmp_17 : _GEN_646; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_652 = cs_100 ? _GEN_650 : _GEN_646; // @[MemMap.scala 164:16]
  wire  _GEN_654 = cs_100 | _GEN_648; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_655 = ~cpu_io_as ? 1'h0 : _GEN_654; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_656 = offset_17 == 24'h4 ? 1'h0 : _GEN_550; // @[Main.scala 222:{26,37}]
  wire  _GEN_658 = cs_18 & readStrobe ? _GEN_656 : _GEN_550; // @[MemMap.scala 180:30]
  wire [15:0] _GEN_660 = cs_18 & readStrobe ? {{13'd0}, _dinReg_T_5} : _GEN_652; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_661 = cs_18 & readStrobe | _GEN_655; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_662 = ~cpu_io_as ? 1'h0 : _GEN_661; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_663 = cs_19 & _upperWriteStrobe_T_3 | _GEN_662; // @[MemMap.scala 154:{27,38}]
  wire  _GEN_664 = ~cpu_io_as ? 1'h0 : _GEN_663; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_665 = cs_20 & writeStrobe | _GEN_557; // @[MemMap.scala 192:31 Main.scala 258:68]
  wire  _GEN_666 = cs_20 & writeStrobe | _GEN_664; // @[MemMap.scala 192:31 194:18]
  wire  _GEN_667 = ~cpu_io_as ? 1'h0 : _GEN_666; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_668 = readStrobe ? 16'h0 : _GEN_660; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_669 = cs_21 ? _GEN_668 : _GEN_660; // @[MemMap.scala 164:16]
  wire  _GEN_670 = cs_21 | _GEN_667; // @[MemMap.scala 164:16 170:18]
  wire  cs_105 = addr_230 >= 24'h800f00 & addr_230 <= 24'h800f03; // @[Util.scala 64:67]
  wire  _GEN_671 = ~cpu_io_as ? 1'h0 : _GEN_670; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_672 = cs_105 & readStrobe ? 16'h0 : _GEN_669; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_673 = cs_105 & readStrobe | _GEN_671; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_674 = ~cpu_io_as ? 1'h0 : _GEN_673; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_675 = cs_22 ? layerRegs_0_io_mem_dout : _GEN_672; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_676 = cs_22 | _GEN_674; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_677 = ~cpu_io_as ? 1'h0 : _GEN_676; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_678 = cs_23 ? layerRegs_1_io_mem_dout : _GEN_675; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_679 = cs_23 | _GEN_677; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_680 = ~cpu_io_as ? 1'h0 : _GEN_679; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_681 = cs_77 ? layerRegs_2_io_mem_dout : _GEN_678; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_682 = cs_77 | _GEN_680; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_683 = ~cpu_io_as ? 1'h0 : _GEN_682; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_684 = cs_78 ? paletteRam_io_portA_dout : _GEN_681; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_685 = cs_78 | _GEN_683; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_686 = ~cpu_io_as ? 1'h0 : _GEN_685; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_687 = cs_211 & readStrobe ? input0 : _GEN_684; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_688 = cs_211 & readStrobe | _GEN_686; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_689 = ~cpu_io_as ? 1'h0 : _GEN_688; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_690 = cs_80 & readStrobe ? input1 : _GEN_687; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_691 = cs_80 & readStrobe | _GEN_689; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_692 = ~cpu_io_as ? 1'h0 : _GEN_691; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_693 = cs_112 & _upperWriteStrobe_T_3 | _GEN_692; // @[MemMap.scala 154:{27,38}]
  wire  _GEN_694 = io_gameIndex == 4'h3 ? _GEN_693 : _GEN_508; // @[Main.scala 326:41]
  wire  _GEN_697 = io_gameIndex == 4'h3 ? cs_2 & readStrobe : _GEN_511; // @[Main.scala 326:41 MemMap.scala 128:14]
  wire [23:0] _GEN_698 = io_gameIndex == 4'h3 ? addr_230 : _GEN_512; // @[Main.scala 326:41 MemMap.scala 129:16]
  wire [15:0] _GEN_699 = io_gameIndex == 4'h3 ? _GEN_690 : _GEN_513; // @[Main.scala 326:41]
  wire  _GEN_700 = io_gameIndex == 4'h3 ? cs_3 & readStrobe : _GEN_514; // @[Main.scala 326:41 MemMap.scala 103:14]
  wire  _GEN_701 = io_gameIndex == 4'h3 ? cs_3 & writeStrobe : _GEN_515; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire [22:0] _GEN_702 = io_gameIndex == 4'h3 ? cpu_io_addr : _GEN_516; // @[Main.scala 326:41 MemMap.scala 105:16]
  wire [1:0] _GEN_703 = io_gameIndex == 4'h3 ? _mainRam_io_mask_T : _GEN_517; // @[Main.scala 326:41 MemMap.scala 106:16]
  wire  _GEN_705 = io_gameIndex == 4'h3 ? cs_4 & readStrobe : _GEN_519; // @[Main.scala 326:41 MemMap.scala 103:14]
  wire  _GEN_706 = io_gameIndex == 4'h3 ? cs_4 & writeStrobe : _GEN_520; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire [22:0] _GEN_707 = io_gameIndex == 4'h3 ? cpu_io_addr : _GEN_521; // @[Main.scala 326:41 MemMap.scala 105:16]
  wire [1:0] _GEN_708 = io_gameIndex == 4'h3 ? _mainRam_io_mask_T : _GEN_522; // @[Main.scala 326:41 MemMap.scala 106:16]
  wire [15:0] _GEN_709 = io_gameIndex == 4'h3 ? cpu_io_dout : _GEN_523; // @[Main.scala 326:41 MemMap.scala 107:15]
  wire  _GEN_710 = io_gameIndex == 4'h3 ? cs_5 & readStrobe : _GEN_524; // @[Main.scala 326:41 MemMap.scala 103:14]
  wire  _GEN_711 = io_gameIndex == 4'h3 ? cs_5 & writeStrobe : _GEN_525; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire  _GEN_713 = io_gameIndex == 4'h3 ? cs_6 & readStrobe : _GEN_527; // @[Main.scala 326:41 MemMap.scala 103:14]
  wire  _GEN_714 = io_gameIndex == 4'h3 ? cs_6 & writeStrobe : _GEN_528; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire  _GEN_716 = io_gameIndex == 4'h3 ? cs_7 & readStrobe : _GEN_530; // @[Main.scala 326:41 MemMap.scala 103:14]
  wire  _GEN_717 = io_gameIndex == 4'h3 ? cs_7 & writeStrobe : _GEN_531; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire  _GEN_719 = io_gameIndex == 4'h3 ? cs_9 & readStrobe : _GEN_533; // @[Main.scala 326:41 MemMap.scala 103:14]
  wire  _GEN_720 = io_gameIndex == 4'h3 ? cs_9 & writeStrobe : _GEN_534; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire  _GEN_722 = io_gameIndex == 4'h3 ? cs_11 & readStrobe : _GEN_536; // @[Main.scala 326:41 MemMap.scala 103:14]
  wire  _GEN_723 = io_gameIndex == 4'h3 ? cs_11 & writeStrobe : _GEN_537; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire  _GEN_725 = io_gameIndex == 4'h3 ? cs_12 & readStrobe : _GEN_539; // @[Main.scala 326:41 MemMap.scala 103:14]
  wire  _GEN_726 = io_gameIndex == 4'h3 ? cs_12 & writeStrobe : _GEN_540; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire  _GEN_728 = io_gameIndex == 4'h3 ? cs_14 & readStrobe : _GEN_542; // @[Main.scala 326:41 MemMap.scala 103:14]
  wire  _GEN_729 = io_gameIndex == 4'h3 ? cs_14 & writeStrobe : _GEN_543; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire  _GEN_731 = io_gameIndex == 4'h3 & (cs_96 & readStrobe); // @[Main.scala 326:41 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_732 = io_gameIndex == 4'h3 & (cs_96 & writeStrobe); // @[Main.scala 326:41 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_736 = io_gameIndex == 4'h3 & (cs_97 & readStrobe); // @[Main.scala 326:41 MemMap.scala 103:14 MemIO.scala 317:8]
  wire  _GEN_737 = io_gameIndex == 4'h3 & (cs_97 & writeStrobe); // @[Main.scala 326:41 MemMap.scala 104:14 MemIO.scala 318:8]
  wire  _GEN_739 = io_gameIndex == 4'h3 ? cs_99 & readStrobe : _GEN_545; // @[Main.scala 326:41 MemMap.scala 103:14]
  wire  _GEN_740 = io_gameIndex == 4'h3 ? cs_99 & writeStrobe : _GEN_546; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire [22:0] _GEN_741 = io_gameIndex == 4'h3 ? cpu_io_addr : {{10'd0}, _GEN_547}; // @[Main.scala 326:41 MemMap.scala 105:16]
  wire  _GEN_744 = io_gameIndex == 4'h3 ? _GEN_658 : _GEN_550; // @[Main.scala 326:41]
  wire  _GEN_747 = io_gameIndex == 4'h3 ? mem_wr : _GEN_553; // @[Main.scala 326:41 MemIO.scala 305:8]
  wire [2:0] _GEN_748 = io_gameIndex == 4'h3 ? mem_addr : _GEN_554; // @[Main.scala 326:41 MemIO.scala 306:10]
  wire [15:0] _GEN_750 = io_gameIndex == 4'h3 ? _GEN_193 : _GEN_556; // @[Main.scala 326:41 MemIO.scala 308:9]
  wire  _GEN_751 = io_gameIndex == 4'h3 ? _GEN_665 : _GEN_557; // @[Main.scala 326:41]
  wire  _GEN_753 = io_gameIndex == 4'h3 ? cs_22 & writeStrobe : _GEN_559; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire  _GEN_756 = io_gameIndex == 4'h3 ? cs_23 & writeStrobe : _GEN_562; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire  _GEN_759 = io_gameIndex == 4'h3 ? cs_77 & writeStrobe : _GEN_565; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire  _GEN_762 = io_gameIndex == 4'h3 ? cs_78 & readStrobe : _GEN_568; // @[Main.scala 326:41 MemMap.scala 103:14]
  wire  _GEN_763 = io_gameIndex == 4'h3 ? cs_78 & writeStrobe : _GEN_569; // @[Main.scala 326:41 MemMap.scala 104:14]
  wire [22:0] _GEN_764 = io_gameIndex == 4'h3 ? cpu_io_addr : _GEN_570; // @[Main.scala 326:41 MemMap.scala 105:16]
  wire  _GEN_768 = ~cpu_io_as ? 1'h0 : _GEN_694; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_769 = cs_2 & cpu_io_rw & io_progRom_valid ? io_progRom_dout : _GEN_699; // @[MemMap.scala 130:39 131:16]
  wire  _GEN_770 = cs_2 & cpu_io_rw & io_progRom_valid | _GEN_768; // @[MemMap.scala 130:39 132:18]
  wire  cs_114 = addr_230 >= 24'h57e & addr_230 <= 24'h581; // @[Util.scala 64:67]
  wire  _GEN_771 = ~cpu_io_as ? 1'h0 : _GEN_770; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_772 = cs_114 & writeStrobe | _GEN_771; // @[MemMap.scala 192:31 194:18]
  wire  _GEN_773 = ~cpu_io_as ? 1'h0 : _GEN_772; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_774 = cs_3 ? mainRam_io_dout : _GEN_769; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_775 = cs_3 | _GEN_773; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_776 = ~cpu_io_as ? 1'h0 : _GEN_775; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_777 = cs_4 ? io_soundCtrl_ymz_dout : _GEN_774; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_778 = cs_4 | _GEN_776; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_779 = ~cpu_io_as ? 1'h0 : _GEN_778; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_780 = cs_5 ? spriteRam_io_portA_dout : _GEN_777; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_781 = cs_5 | _GEN_779; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_782 = ~cpu_io_as ? 1'h0 : _GEN_781; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_783 = cs_6 ? vram16x16_0_io_portA_dout : _GEN_780; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_784 = cs_6 | _GEN_782; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_785 = ~cpu_io_as ? 1'h0 : _GEN_784; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_786 = cs_7 ? lineRam_0_io_portA_dout : _GEN_783; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_787 = cs_7 | _GEN_785; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_788 = ~cpu_io_as ? 1'h0 : _GEN_787; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_18; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_790 = readStrobe ? tmp_18 : _GEN_786; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_792 = cs_8 ? _GEN_790 : _GEN_786; // @[MemMap.scala 164:16]
  wire  _GEN_794 = cs_8 | _GEN_788; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_795 = ~cpu_io_as ? 1'h0 : _GEN_794; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_796 = cs_9 ? vram8x8_0_io_portA_dout : _GEN_792; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_797 = cs_9 | _GEN_795; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_798 = ~cpu_io_as ? 1'h0 : _GEN_797; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_19; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_800 = readStrobe ? tmp_19 : _GEN_796; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_802 = cs_10 ? _GEN_800 : _GEN_796; // @[MemMap.scala 164:16]
  wire  _GEN_804 = cs_10 | _GEN_798; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_805 = ~cpu_io_as ? 1'h0 : _GEN_804; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_806 = cs_11 ? vram16x16_1_io_portA_dout : _GEN_802; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_807 = cs_11 | _GEN_805; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_808 = ~cpu_io_as ? 1'h0 : _GEN_807; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_809 = cs_12 ? lineRam_1_io_portA_dout : _GEN_806; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_810 = cs_12 | _GEN_808; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_811 = ~cpu_io_as ? 1'h0 : _GEN_810; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_20; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_813 = readStrobe ? tmp_20 : _GEN_809; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_815 = cs_13 ? _GEN_813 : _GEN_809; // @[MemMap.scala 164:16]
  wire  _GEN_817 = cs_13 | _GEN_811; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_818 = ~cpu_io_as ? 1'h0 : _GEN_817; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_819 = cs_14 ? vram8x8_1_io_portA_dout : _GEN_815; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_820 = cs_14 | _GEN_818; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_821 = ~cpu_io_as ? 1'h0 : _GEN_820; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_21; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_823 = readStrobe ? tmp_21 : _GEN_819; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_825 = cs_15 ? _GEN_823 : _GEN_819; // @[MemMap.scala 164:16]
  wire  _GEN_827 = cs_15 | _GEN_821; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_828 = ~cpu_io_as ? 1'h0 : _GEN_827; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_829 = cs_96 ? vram16x16_2_io_portA_dout : _GEN_825; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_830 = cs_96 | _GEN_828; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_831 = ~cpu_io_as ? 1'h0 : _GEN_830; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_832 = cs_97 ? lineRam_2_io_portA_dout : _GEN_829; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_833 = cs_97 | _GEN_831; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_834 = ~cpu_io_as ? 1'h0 : _GEN_833; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_22; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_836 = readStrobe ? tmp_22 : _GEN_832; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_838 = cs_98 ? _GEN_836 : _GEN_832; // @[MemMap.scala 164:16]
  wire  _GEN_840 = cs_98 | _GEN_834; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_841 = ~cpu_io_as ? 1'h0 : _GEN_840; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_842 = cs_99 ? vram8x8_2_io_portA_dout : _GEN_838; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_843 = cs_99 | _GEN_841; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_844 = ~cpu_io_as ? 1'h0 : _GEN_843; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_23; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_846 = readStrobe ? tmp_23 : _GEN_842; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_848 = cs_100 ? _GEN_846 : _GEN_842; // @[MemMap.scala 164:16]
  wire  _GEN_850 = cs_100 | _GEN_844; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_851 = ~cpu_io_as ? 1'h0 : _GEN_850; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_852 = offset_17 == 24'h4 ? 1'h0 : _GEN_744; // @[Main.scala 222:{26,37}]
  wire  _GEN_854 = cs_18 & readStrobe ? _GEN_852 : _GEN_744; // @[MemMap.scala 180:30]
  wire [15:0] _GEN_856 = cs_18 & readStrobe ? {{13'd0}, _dinReg_T_5} : _GEN_848; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_857 = cs_18 & readStrobe | _GEN_851; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_858 = ~cpu_io_as ? 1'h0 : _GEN_857; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_859 = cs_19 & _upperWriteStrobe_T_3 | _GEN_858; // @[MemMap.scala 154:{27,38}]
  wire  _GEN_860 = ~cpu_io_as ? 1'h0 : _GEN_859; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_861 = cs_20 & writeStrobe | _GEN_751; // @[MemMap.scala 192:31 Main.scala 258:68]
  wire  _GEN_862 = cs_20 & writeStrobe | _GEN_860; // @[MemMap.scala 192:31 194:18]
  wire  _GEN_863 = ~cpu_io_as ? 1'h0 : _GEN_862; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_864 = readStrobe ? 16'h0 : _GEN_856; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_865 = cs_21 ? _GEN_864 : _GEN_856; // @[MemMap.scala 164:16]
  wire  _GEN_866 = cs_21 | _GEN_863; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_867 = ~cpu_io_as ? 1'h0 : _GEN_866; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_868 = cs_22 ? layerRegs_0_io_mem_dout : _GEN_865; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_869 = cs_22 | _GEN_867; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_870 = ~cpu_io_as ? 1'h0 : _GEN_869; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_871 = cs_23 ? layerRegs_1_io_mem_dout : _GEN_868; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_872 = cs_23 | _GEN_870; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_873 = ~cpu_io_as ? 1'h0 : _GEN_872; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_874 = cs_77 ? layerRegs_2_io_mem_dout : _GEN_871; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_875 = cs_77 | _GEN_873; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_876 = ~cpu_io_as ? 1'h0 : _GEN_875; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_877 = cs_78 ? paletteRam_io_portA_dout : _GEN_874; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_878 = cs_78 | _GEN_876; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_879 = ~cpu_io_as ? 1'h0 : _GEN_878; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_880 = cs_179 & readStrobe ? input0 : _GEN_877; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_881 = cs_179 & readStrobe | _GEN_879; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_882 = ~cpu_io_as ? 1'h0 : _GEN_881; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_883 = _eepromMem_wr_T_4 | _GEN_882; // @[MemMap.scala 192:31 194:18]
  wire  cs_143 = addr_230 >= 24'hd00012 & addr_230 <= 24'hd00012; // @[Util.scala 64:67]
  wire  _GEN_884 = ~cpu_io_as ? 1'h0 : _GEN_883; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_885 = cs_143 & readStrobe ? input1 : _GEN_880; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_886 = cs_143 & readStrobe | _GEN_884; // @[MemMap.scala 180:30 182:18]
  wire  cs_144 = addr_230 >= 24'hd00014 & addr_230 <= 24'hd00014; // @[Util.scala 64:67]
  wire  _GEN_887 = ~cpu_io_as ? 1'h0 : _GEN_886; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_888 = cs_144 & readStrobe ? io_dips_0 : _GEN_885; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_889 = cs_144 & readStrobe | _GEN_887; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_890 = ~cpu_io_as ? 1'h0 : _GEN_889; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_891 = cs_144 & writeStrobe | _GEN_890; // @[MemMap.scala 192:31 194:18]
  wire  _GEN_892 = io_gameIndex == 4'h6 ? _GEN_891 : _GEN_694; // @[Main.scala 346:38]
  wire  _GEN_895 = io_gameIndex == 4'h6 ? cs_2 & readStrobe : _GEN_697; // @[Main.scala 346:38 MemMap.scala 128:14]
  wire [23:0] _GEN_896 = io_gameIndex == 4'h6 ? addr_230 : _GEN_698; // @[Main.scala 346:38 MemMap.scala 129:16]
  wire [15:0] _GEN_897 = io_gameIndex == 4'h6 ? _GEN_888 : _GEN_699; // @[Main.scala 346:38]
  wire  _GEN_898 = io_gameIndex == 4'h6 ? cs_3 & readStrobe : _GEN_700; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_899 = io_gameIndex == 4'h6 ? cs_3 & writeStrobe : _GEN_701; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire [22:0] _GEN_900 = io_gameIndex == 4'h6 ? cpu_io_addr : _GEN_702; // @[Main.scala 346:38 MemMap.scala 105:16]
  wire [1:0] _GEN_901 = io_gameIndex == 4'h6 ? _mainRam_io_mask_T : _GEN_703; // @[Main.scala 346:38 MemMap.scala 106:16]
  wire [15:0] _GEN_902 = io_gameIndex == 4'h6 ? cpu_io_dout : _GEN_704; // @[Main.scala 346:38 MemMap.scala 107:15]
  wire  _GEN_903 = io_gameIndex == 4'h6 ? cs_4 & readStrobe : _GEN_705; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_904 = io_gameIndex == 4'h6 ? cs_4 & writeStrobe : _GEN_706; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire [22:0] _GEN_905 = io_gameIndex == 4'h6 ? cpu_io_addr : _GEN_707; // @[Main.scala 346:38 MemMap.scala 105:16]
  wire [1:0] _GEN_906 = io_gameIndex == 4'h6 ? _mainRam_io_mask_T : _GEN_708; // @[Main.scala 346:38 MemMap.scala 106:16]
  wire [15:0] _GEN_907 = io_gameIndex == 4'h6 ? cpu_io_dout : _GEN_709; // @[Main.scala 346:38 MemMap.scala 107:15]
  wire  _GEN_908 = io_gameIndex == 4'h6 ? cs_5 & readStrobe : _GEN_710; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_909 = io_gameIndex == 4'h6 ? cs_5 & writeStrobe : _GEN_711; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire  _GEN_911 = io_gameIndex == 4'h6 ? cs_6 & readStrobe : _GEN_713; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_912 = io_gameIndex == 4'h6 ? cs_6 & writeStrobe : _GEN_714; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire  _GEN_914 = io_gameIndex == 4'h6 ? cs_7 & readStrobe : _GEN_716; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_915 = io_gameIndex == 4'h6 ? cs_7 & writeStrobe : _GEN_717; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire  _GEN_917 = io_gameIndex == 4'h6 ? cs_9 & readStrobe : _GEN_719; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_918 = io_gameIndex == 4'h6 ? cs_9 & writeStrobe : _GEN_720; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire  _GEN_920 = io_gameIndex == 4'h6 ? cs_11 & readStrobe : _GEN_722; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_921 = io_gameIndex == 4'h6 ? cs_11 & writeStrobe : _GEN_723; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire  _GEN_923 = io_gameIndex == 4'h6 ? cs_12 & readStrobe : _GEN_725; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_924 = io_gameIndex == 4'h6 ? cs_12 & writeStrobe : _GEN_726; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire  _GEN_926 = io_gameIndex == 4'h6 ? cs_14 & readStrobe : _GEN_728; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_927 = io_gameIndex == 4'h6 ? cs_14 & writeStrobe : _GEN_729; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire  _GEN_929 = io_gameIndex == 4'h6 ? cs_96 & readStrobe : _GEN_731; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_930 = io_gameIndex == 4'h6 ? cs_96 & writeStrobe : _GEN_732; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire [22:0] _GEN_931 = io_gameIndex == 4'h6 ? cpu_io_addr : _GEN_191; // @[Main.scala 346:38 MemMap.scala 105:16]
  wire [1:0] _GEN_932 = io_gameIndex == 4'h6 ? _mainRam_io_mask_T : _mainRam_io_mask_T; // @[Main.scala 346:38 MemMap.scala 106:16]
  wire [15:0] _GEN_933 = io_gameIndex == 4'h6 ? cpu_io_dout : _GEN_193; // @[Main.scala 346:38 MemMap.scala 107:15]
  wire  _GEN_934 = io_gameIndex == 4'h6 ? cs_97 & readStrobe : _GEN_736; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_935 = io_gameIndex == 4'h6 ? cs_97 & writeStrobe : _GEN_737; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire  _GEN_937 = io_gameIndex == 4'h6 ? cs_99 & readStrobe : _GEN_739; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_938 = io_gameIndex == 4'h6 ? cs_99 & writeStrobe : _GEN_740; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire [22:0] _GEN_939 = io_gameIndex == 4'h6 ? cpu_io_addr : _GEN_741; // @[Main.scala 346:38 MemMap.scala 105:16]
  wire  _GEN_942 = io_gameIndex == 4'h6 ? _GEN_854 : _GEN_744; // @[Main.scala 346:38]
  wire  _GEN_945 = io_gameIndex == 4'h6 ? mem_wr : _GEN_747; // @[Main.scala 346:38 MemIO.scala 305:8]
  wire [2:0] _GEN_946 = io_gameIndex == 4'h6 ? mem_addr : _GEN_748; // @[Main.scala 346:38 MemIO.scala 306:10]
  wire [15:0] _GEN_948 = io_gameIndex == 4'h6 ? _GEN_193 : _GEN_750; // @[Main.scala 346:38 MemIO.scala 308:9]
  wire  _GEN_949 = io_gameIndex == 4'h6 ? _GEN_861 : _GEN_751; // @[Main.scala 346:38]
  wire  _GEN_951 = io_gameIndex == 4'h6 ? cs_22 & writeStrobe : _GEN_753; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire  _GEN_954 = io_gameIndex == 4'h6 ? cs_23 & writeStrobe : _GEN_756; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire  _GEN_957 = io_gameIndex == 4'h6 ? cs_77 & writeStrobe : _GEN_759; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire  _GEN_960 = io_gameIndex == 4'h6 ? cs_78 & readStrobe : _GEN_762; // @[Main.scala 346:38 MemMap.scala 103:14]
  wire  _GEN_961 = io_gameIndex == 4'h6 ? cs_78 & writeStrobe : _GEN_763; // @[Main.scala 346:38 MemMap.scala 104:14]
  wire [22:0] _GEN_962 = io_gameIndex == 4'h6 ? cpu_io_addr : _GEN_764; // @[Main.scala 346:38 MemMap.scala 105:16]
  wire  _GEN_964 = ~cpu_io_as ? 1'h0 : _GEN_892; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_965 = cs_2 & cpu_io_rw & io_progRom_valid ? io_progRom_dout : _GEN_897; // @[MemMap.scala 130:39 131:16]
  wire  _GEN_966 = cs_2 & cpu_io_rw & io_progRom_valid | _GEN_964; // @[MemMap.scala 130:39 132:18]
  wire  cs_147 = addr_230 >= 24'h200000 & addr_230 <= 24'h20ffff; // @[Util.scala 64:67]
  wire  _GEN_967 = ~cpu_io_as ? 1'h0 : _GEN_966; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_968 = cs_147 ? mainRam_io_dout : _GEN_965; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_969 = cs_147 | _GEN_967; // @[MemMap.scala 108:16 110:18]
  wire  cs_148 = addr_230 >= 24'h210000 & addr_230 <= 24'h2fffff; // @[Util.scala 64:67]
  wire  _GEN_970 = ~cpu_io_as ? 1'h0 : _GEN_969; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_971 = cs_148 & readStrobe ? 16'h0 : _GEN_968; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_972 = cs_148 & readStrobe | _GEN_970; // @[MemMap.scala 180:30 182:18]
  wire  cs_149 = addr_230 >= 24'h300000 & addr_230 <= 24'h300007; // @[Util.scala 64:67]
  wire  _GEN_973 = ~cpu_io_as ? 1'h0 : _GEN_972; // @[MemMap.scala 226:{19,30}]
  wire  dinReg_a_5 = offset_3 == 24'h0 & agalletIrq; // @[Main.scala 219:28]
  wire  _GEN_974 = offset_3 == 24'h4 ? 1'h0 : _GEN_942; // @[Main.scala 222:{26,37}]
  wire  _dinReg_T_32 = ~dinReg_a_5; // @[Main.scala 224:9]
  wire [2:0] _dinReg_T_35 = {_dinReg_T_32,1'h1,_dinReg_T_4}; // @[Cat.scala 33:92]
  wire  _GEN_976 = cs_149 & readStrobe ? _GEN_974 : _GEN_942; // @[MemMap.scala 180:30]
  wire [15:0] _GEN_978 = cs_149 & readStrobe ? {{13'd0}, _dinReg_T_35} : _GEN_971; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_979 = cs_149 & readStrobe | _GEN_973; // @[MemMap.scala 180:30 182:18]
  wire  cs_150 = addr_230 >= 24'h300000 & addr_230 <= 24'h30000f; // @[Util.scala 64:67]
  wire  _GEN_980 = ~cpu_io_as ? 1'h0 : _GEN_979; // @[MemMap.scala 226:{19,30}]
  wire  mem_5_wr = cs_150 & writeStrobe; // @[MemMap.scala 150:20]
  wire  _GEN_981 = cs_150 & _upperWriteStrobe_T_3 | _GEN_980; // @[MemMap.scala 154:{27,38}]
  wire  cs_151 = addr_230 >= 24'h300008 & addr_230 <= 24'h300008; // @[Util.scala 64:67]
  wire  _GEN_982 = ~cpu_io_as ? 1'h0 : _GEN_981; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_983 = cs_151 & writeStrobe | _GEN_949; // @[MemMap.scala 192:31 Main.scala 258:68]
  wire  _GEN_984 = cs_151 & writeStrobe | _GEN_982; // @[MemMap.scala 192:31 194:18]
  wire  cs_152 = addr_230 >= 24'h30000a & addr_230 <= 24'h30007f; // @[Util.scala 64:67]
  wire  _GEN_985 = ~cpu_io_as ? 1'h0 : _GEN_984; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_986 = readStrobe ? 16'h0 : _GEN_978; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_987 = cs_152 ? _GEN_986 : _GEN_978; // @[MemMap.scala 164:16]
  wire  _GEN_988 = cs_152 | _GEN_985; // @[MemMap.scala 164:16 170:18]
  wire  cs_153 = addr_230 >= 24'h300080 & addr_230 <= 24'h3fffff; // @[Util.scala 64:67]
  wire  _GEN_989 = ~cpu_io_as ? 1'h0 : _GEN_988; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_990 = cs_153 & readStrobe ? 16'h0 : _GEN_987; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_991 = cs_153 & readStrobe | _GEN_989; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_992 = ~cpu_io_as ? 1'h0 : _GEN_991; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_993 = cs_5 ? spriteRam_io_portA_dout : _GEN_990; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_994 = cs_5 | _GEN_992; // @[MemMap.scala 108:16 110:18]
  wire  cs_155 = addr_230 >= 24'h410000 & addr_230 <= 24'h4fffff; // @[Util.scala 64:67]
  wire  _GEN_995 = ~cpu_io_as ? 1'h0 : _GEN_994; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_996 = cs_155 & readStrobe ? 16'h0 : _GEN_993; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_997 = cs_155 & readStrobe | _GEN_995; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_998 = ~cpu_io_as ? 1'h0 : _GEN_997; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_999 = cs_6 ? vram16x16_0_io_portA_dout : _GEN_996; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1000 = cs_6 | _GEN_998; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1001 = ~cpu_io_as ? 1'h0 : _GEN_1000; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1002 = cs_7 ? lineRam_0_io_portA_dout : _GEN_999; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1003 = cs_7 | _GEN_1001; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1004 = ~cpu_io_as ? 1'h0 : _GEN_1003; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_24; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1006 = readStrobe ? tmp_24 : _GEN_1002; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1008 = cs_8 ? _GEN_1006 : _GEN_1002; // @[MemMap.scala 164:16]
  wire  _GEN_1010 = cs_8 | _GEN_1004; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_1011 = ~cpu_io_as ? 1'h0 : _GEN_1010; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1012 = cs_9 ? vram8x8_0_io_portA_dout : _GEN_1008; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1013 = cs_9 | _GEN_1011; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1014 = ~cpu_io_as ? 1'h0 : _GEN_1013; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_25; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1016 = readStrobe ? tmp_25 : _GEN_1012; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1018 = cs_10 ? _GEN_1016 : _GEN_1012; // @[MemMap.scala 164:16]
  wire  _GEN_1020 = cs_10 | _GEN_1014; // @[MemMap.scala 164:16 170:18]
  wire  cs_161 = addr_230 >= 24'h508000 & addr_230 <= 24'h5fffff; // @[Util.scala 64:67]
  wire  _GEN_1021 = ~cpu_io_as ? 1'h0 : _GEN_1020; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1022 = cs_161 & readStrobe ? 16'h0 : _GEN_1018; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_1023 = cs_161 & readStrobe | _GEN_1021; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_1024 = ~cpu_io_as ? 1'h0 : _GEN_1023; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1025 = cs_11 ? vram16x16_1_io_portA_dout : _GEN_1022; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1026 = cs_11 | _GEN_1024; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1027 = ~cpu_io_as ? 1'h0 : _GEN_1026; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1028 = cs_12 ? lineRam_1_io_portA_dout : _GEN_1025; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1029 = cs_12 | _GEN_1027; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1030 = ~cpu_io_as ? 1'h0 : _GEN_1029; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_26; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1032 = readStrobe ? tmp_26 : _GEN_1028; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1034 = cs_13 ? _GEN_1032 : _GEN_1028; // @[MemMap.scala 164:16]
  wire  _GEN_1036 = cs_13 | _GEN_1030; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_1037 = ~cpu_io_as ? 1'h0 : _GEN_1036; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1038 = cs_14 ? vram8x8_1_io_portA_dout : _GEN_1034; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1039 = cs_14 | _GEN_1037; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1040 = ~cpu_io_as ? 1'h0 : _GEN_1039; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_27; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1042 = readStrobe ? tmp_27 : _GEN_1038; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1044 = cs_15 ? _GEN_1042 : _GEN_1038; // @[MemMap.scala 164:16]
  wire  _GEN_1046 = cs_15 | _GEN_1040; // @[MemMap.scala 164:16 170:18]
  wire  cs_167 = addr_230 >= 24'h608000 & addr_230 <= 24'h6fffff; // @[Util.scala 64:67]
  wire  _GEN_1047 = ~cpu_io_as ? 1'h0 : _GEN_1046; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1048 = cs_167 & readStrobe ? 16'h0 : _GEN_1044; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_1049 = cs_167 & readStrobe | _GEN_1047; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_1050 = ~cpu_io_as ? 1'h0 : _GEN_1049; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1051 = cs_96 ? vram16x16_2_io_portA_dout : _GEN_1048; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1052 = cs_96 | _GEN_1050; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1053 = ~cpu_io_as ? 1'h0 : _GEN_1052; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1054 = cs_97 ? lineRam_2_io_portA_dout : _GEN_1051; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1055 = cs_97 | _GEN_1053; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1056 = ~cpu_io_as ? 1'h0 : _GEN_1055; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_28; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1058 = readStrobe ? tmp_28 : _GEN_1054; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1060 = cs_98 ? _GEN_1058 : _GEN_1054; // @[MemMap.scala 164:16]
  wire  _GEN_1062 = cs_98 | _GEN_1056; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_1063 = ~cpu_io_as ? 1'h0 : _GEN_1062; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1064 = cs_99 ? vram8x8_2_io_portA_dout : _GEN_1060; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1065 = cs_99 | _GEN_1063; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1066 = ~cpu_io_as ? 1'h0 : _GEN_1065; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_29; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1068 = readStrobe ? tmp_29 : _GEN_1064; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1070 = cs_100 ? _GEN_1068 : _GEN_1064; // @[MemMap.scala 164:16]
  wire  _GEN_1072 = cs_100 | _GEN_1066; // @[MemMap.scala 164:16 170:18]
  wire  cs_173 = addr_230 >= 24'h800000 & addr_230 <= 24'h800003; // @[Util.scala 64:67]
  wire  _GEN_1073 = ~cpu_io_as ? 1'h0 : _GEN_1072; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1074 = cs_173 ? io_soundCtrl_ymz_dout : _GEN_1070; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1075 = cs_173 | _GEN_1073; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1076 = ~cpu_io_as ? 1'h0 : _GEN_1075; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1077 = cs_22 ? layerRegs_0_io_mem_dout : _GEN_1074; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1078 = cs_22 | _GEN_1076; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1079 = ~cpu_io_as ? 1'h0 : _GEN_1078; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1080 = cs_23 ? layerRegs_1_io_mem_dout : _GEN_1077; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1081 = cs_23 | _GEN_1079; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1082 = ~cpu_io_as ? 1'h0 : _GEN_1081; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1083 = cs_77 ? layerRegs_2_io_mem_dout : _GEN_1080; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1084 = cs_77 | _GEN_1082; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1085 = ~cpu_io_as ? 1'h0 : _GEN_1084; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1086 = cs_78 ? paletteRam_io_portA_dout : _GEN_1083; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1087 = cs_78 | _GEN_1085; // @[MemMap.scala 108:16 110:18]
  wire  cs_178 = addr_230 >= 24'hd00010 & addr_230 <= 24'hd00014; // @[Util.scala 64:67]
  wire  _GEN_1088 = ~cpu_io_as ? 1'h0 : _GEN_1087; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1089 = readStrobe ? 16'h0 : _GEN_1086; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1090 = cs_178 ? _GEN_1089 : _GEN_1086; // @[MemMap.scala 164:16]
  wire  _GEN_1091 = cs_178 | _GEN_1088; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_1092 = ~cpu_io_as ? 1'h0 : _GEN_1091; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_1093 = cs_179 & _upperWriteStrobe_T_3 | _GEN_1092; // @[MemMap.scala 154:{27,38}]
  wire  _GEN_1094 = ~cpu_io_as ? 1'h0 : _GEN_1093; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1095 = cs_179 & readStrobe ? input0 : _GEN_1090; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_1096 = cs_179 & readStrobe | _GEN_1094; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_1097 = ~cpu_io_as ? 1'h0 : _GEN_1096; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1098 = cs_143 & readStrobe ? input1 : _GEN_1095; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_1099 = cs_143 & readStrobe | _GEN_1097; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_1100 = _cs_T ? _GEN_1099 : _GEN_892; // @[Main.scala 368:41]
  wire  _GEN_1103 = _cs_T ? cs_2 & readStrobe : _GEN_895; // @[Main.scala 368:41 MemMap.scala 128:14]
  wire [23:0] _GEN_1104 = _cs_T ? addr_230 : _GEN_896; // @[Main.scala 368:41 MemMap.scala 129:16]
  wire [15:0] _GEN_1105 = _cs_T ? _GEN_1098 : _GEN_897; // @[Main.scala 368:41]
  wire  _GEN_1106 = _cs_T ? cs_147 & readStrobe : _GEN_898; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1107 = _cs_T ? cs_147 & writeStrobe : _GEN_899; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire [22:0] _GEN_1108 = _cs_T ? cpu_io_addr : _GEN_900; // @[Main.scala 368:41 MemMap.scala 105:16]
  wire [1:0] _GEN_1109 = _cs_T ? _mainRam_io_mask_T : _GEN_901; // @[Main.scala 368:41 MemMap.scala 106:16]
  wire [15:0] _GEN_1110 = _cs_T ? cpu_io_dout : _GEN_902; // @[Main.scala 368:41 MemMap.scala 107:15]
  wire  _GEN_1111 = _cs_T ? _GEN_976 : _GEN_942; // @[Main.scala 368:41]
  wire  _GEN_1114 = _cs_T ? mem_5_wr : _GEN_945; // @[Main.scala 368:41 MemIO.scala 305:8]
  wire [2:0] _GEN_1115 = _cs_T ? mem_addr : _GEN_946; // @[Main.scala 368:41 MemIO.scala 306:10]
  wire [15:0] _GEN_1117 = _cs_T ? _GEN_193 : _GEN_948; // @[Main.scala 368:41 MemIO.scala 308:9]
  wire  _GEN_1118 = _cs_T ? _GEN_983 : _GEN_949; // @[Main.scala 368:41]
  wire  _GEN_1119 = _cs_T ? cs_5 & readStrobe : _GEN_908; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1120 = _cs_T ? cs_5 & writeStrobe : _GEN_909; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire  _GEN_1122 = _cs_T ? cs_6 & readStrobe : _GEN_911; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1123 = _cs_T ? cs_6 & writeStrobe : _GEN_912; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire  _GEN_1125 = _cs_T ? cs_7 & readStrobe : _GEN_914; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1126 = _cs_T ? cs_7 & writeStrobe : _GEN_915; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire  _GEN_1128 = _cs_T ? cs_9 & readStrobe : _GEN_917; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1129 = _cs_T ? cs_9 & writeStrobe : _GEN_918; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire  _GEN_1131 = _cs_T ? cs_11 & readStrobe : _GEN_920; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1132 = _cs_T ? cs_11 & writeStrobe : _GEN_921; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire  _GEN_1134 = _cs_T ? cs_12 & readStrobe : _GEN_923; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1135 = _cs_T ? cs_12 & writeStrobe : _GEN_924; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire  _GEN_1137 = _cs_T ? cs_14 & readStrobe : _GEN_926; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1138 = _cs_T ? cs_14 & writeStrobe : _GEN_927; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire  _GEN_1140 = _cs_T ? cs_96 & readStrobe : _GEN_929; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1141 = _cs_T ? cs_96 & writeStrobe : _GEN_930; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire [22:0] _GEN_1142 = _cs_T ? cpu_io_addr : _GEN_931; // @[Main.scala 368:41 MemMap.scala 105:16]
  wire [1:0] _GEN_1143 = _cs_T ? _mainRam_io_mask_T : _GEN_932; // @[Main.scala 368:41 MemMap.scala 106:16]
  wire [15:0] _GEN_1144 = _cs_T ? cpu_io_dout : _GEN_933; // @[Main.scala 368:41 MemMap.scala 107:15]
  wire  _GEN_1145 = _cs_T ? cs_97 & readStrobe : _GEN_934; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1146 = _cs_T ? cs_97 & writeStrobe : _GEN_935; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire  _GEN_1148 = _cs_T ? cs_99 & readStrobe : _GEN_937; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1149 = _cs_T ? cs_99 & writeStrobe : _GEN_938; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire [22:0] _GEN_1150 = _cs_T ? cpu_io_addr : _GEN_939; // @[Main.scala 368:41 MemMap.scala 105:16]
  wire [1:0] _GEN_1151 = _cs_T ? _mainRam_io_mask_T : _GEN_906; // @[Main.scala 368:41 MemMap.scala 106:16]
  wire [15:0] _GEN_1152 = _cs_T ? cpu_io_dout : _GEN_907; // @[Main.scala 368:41 MemMap.scala 107:15]
  wire  _GEN_1153 = _cs_T ? cs_173 & readStrobe : _GEN_903; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1154 = _cs_T ? cs_173 & writeStrobe : _GEN_904; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire [22:0] _GEN_1155 = _cs_T ? cpu_io_addr : _GEN_905; // @[Main.scala 368:41 MemMap.scala 105:16]
  wire  _GEN_1159 = _cs_T ? cs_22 & writeStrobe : _GEN_951; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire  _GEN_1162 = _cs_T ? cs_23 & writeStrobe : _GEN_954; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire  _GEN_1165 = _cs_T ? cs_77 & writeStrobe : _GEN_957; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire  _GEN_1168 = _cs_T ? cs_78 & readStrobe : _GEN_960; // @[Main.scala 368:41 MemMap.scala 103:14]
  wire  _GEN_1169 = _cs_T ? cs_78 & writeStrobe : _GEN_961; // @[Main.scala 368:41 MemMap.scala 104:14]
  wire [22:0] _GEN_1170 = _cs_T ? cpu_io_addr : _GEN_962; // @[Main.scala 368:41 MemMap.scala 105:16]
  wire  _GEN_1176 = ~cpu_io_as ? 1'h0 : _GEN_1100; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1177 = cs_2 & cpu_io_rw & io_progRom_valid ? io_progRom_dout : _GEN_1105; // @[MemMap.scala 130:39 131:16]
  wire  _GEN_1178 = cs_2 & cpu_io_rw & io_progRom_valid | _GEN_1176; // @[MemMap.scala 130:39 132:18]
  wire  cs_183 = addr_230 >= 24'h300000 & addr_230 <= 24'h30ffff; // @[Util.scala 64:67]
  wire  _GEN_1179 = ~cpu_io_as ? 1'h0 : _GEN_1178; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1180 = cs_183 ? mainRam_io_dout : _GEN_1177; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1181 = cs_183 | _GEN_1179; // @[MemMap.scala 108:16 110:18]
  wire  cs_184 = addr_230 >= 24'h408000 & addr_230 <= 24'h408fff; // @[Util.scala 64:67]
  wire  _GEN_1182 = ~cpu_io_as ? 1'h0 : _GEN_1181; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1183 = cs_184 ? paletteRam_io_portA_dout : _GEN_1180; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1184 = cs_184 | _GEN_1182; // @[MemMap.scala 108:16 110:18]
  wire  cs_185 = addr_230 >= 24'h600000 & addr_230 <= 24'h600000; // @[Util.scala 64:67]
  wire  _GEN_1185 = ~cpu_io_as ? 1'h0 : _GEN_1184; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1186 = cs_185 & readStrobe ? 16'h0 : _GEN_1183; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_1187 = cs_185 & readStrobe | _GEN_1185; // @[MemMap.scala 180:30 182:18]
  wire  cs_186 = addr_230 >= 24'h880000 & addr_230 <= 24'h880fff; // @[Util.scala 64:67]
  wire  _GEN_1188 = ~cpu_io_as ? 1'h0 : _GEN_1187; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1189 = cs_186 ? vram16x16_0_io_portA_dout : _GEN_1186; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1190 = cs_186 | _GEN_1188; // @[MemMap.scala 108:16 110:18]
  wire  cs_187 = addr_230 >= 24'h881000 & addr_230 <= 24'h8817ff; // @[Util.scala 64:67]
  wire  _GEN_1191 = ~cpu_io_as ? 1'h0 : _GEN_1190; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1192 = cs_187 ? lineRam_0_io_portA_dout : _GEN_1189; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1193 = cs_187 | _GEN_1191; // @[MemMap.scala 108:16 110:18]
  wire  cs_188 = addr_230 >= 24'h881800 & addr_230 <= 24'h883fff; // @[Util.scala 64:67]
  wire  _GEN_1194 = ~cpu_io_as ? 1'h0 : _GEN_1193; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_30; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1196 = readStrobe ? tmp_30 : _GEN_1192; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1198 = cs_188 ? _GEN_1196 : _GEN_1192; // @[MemMap.scala 164:16]
  wire  _GEN_1200 = cs_188 | _GEN_1194; // @[MemMap.scala 164:16 170:18]
  wire  cs_189 = addr_230 >= 24'h884000 & addr_230 <= 24'h887fff; // @[Util.scala 64:67]
  wire  _GEN_1201 = ~cpu_io_as ? 1'h0 : _GEN_1200; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1202 = cs_189 ? vram8x8_0_io_portA_dout : _GEN_1198; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1203 = cs_189 | _GEN_1201; // @[MemMap.scala 108:16 110:18]
  wire  cs_190 = addr_230 >= 24'h888000 & addr_230 <= 24'h88ffff; // @[Util.scala 64:67]
  wire  _GEN_1204 = ~cpu_io_as ? 1'h0 : _GEN_1203; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_31; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1206 = readStrobe ? tmp_31 : _GEN_1202; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1208 = cs_190 ? _GEN_1206 : _GEN_1202; // @[MemMap.scala 164:16]
  wire  _GEN_1210 = cs_190 | _GEN_1204; // @[MemMap.scala 164:16 170:18]
  wire  cs_191 = addr_230 >= 24'h900000 & addr_230 <= 24'h900fff; // @[Util.scala 64:67]
  wire  _GEN_1211 = ~cpu_io_as ? 1'h0 : _GEN_1210; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1212 = cs_191 ? vram16x16_1_io_portA_dout : _GEN_1208; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1213 = cs_191 | _GEN_1211; // @[MemMap.scala 108:16 110:18]
  wire  cs_192 = addr_230 >= 24'h901000 & addr_230 <= 24'h9017ff; // @[Util.scala 64:67]
  wire  _GEN_1214 = ~cpu_io_as ? 1'h0 : _GEN_1213; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1215 = cs_192 ? lineRam_1_io_portA_dout : _GEN_1212; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1216 = cs_192 | _GEN_1214; // @[MemMap.scala 108:16 110:18]
  wire  cs_193 = addr_230 >= 24'h901800 & addr_230 <= 24'h903fff; // @[Util.scala 64:67]
  wire  _GEN_1217 = ~cpu_io_as ? 1'h0 : _GEN_1216; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_32; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1219 = readStrobe ? tmp_32 : _GEN_1215; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1221 = cs_193 ? _GEN_1219 : _GEN_1215; // @[MemMap.scala 164:16]
  wire  _GEN_1223 = cs_193 | _GEN_1217; // @[MemMap.scala 164:16 170:18]
  wire  cs_194 = addr_230 >= 24'h904000 & addr_230 <= 24'h907fff; // @[Util.scala 64:67]
  wire  _GEN_1224 = ~cpu_io_as ? 1'h0 : _GEN_1223; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1225 = cs_194 ? vram8x8_1_io_portA_dout : _GEN_1221; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1226 = cs_194 | _GEN_1224; // @[MemMap.scala 108:16 110:18]
  wire  cs_195 = addr_230 >= 24'h908000 & addr_230 <= 24'h90ffff; // @[Util.scala 64:67]
  wire  _GEN_1227 = ~cpu_io_as ? 1'h0 : _GEN_1226; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_33; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1229 = readStrobe ? tmp_33 : _GEN_1225; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1231 = cs_195 ? _GEN_1229 : _GEN_1225; // @[MemMap.scala 164:16]
  wire  _GEN_1233 = cs_195 | _GEN_1227; // @[MemMap.scala 164:16 170:18]
  wire  cs_196 = addr_230 >= 24'h980000 & addr_230 <= 24'h980fff; // @[Util.scala 64:67]
  wire  _GEN_1234 = ~cpu_io_as ? 1'h0 : _GEN_1233; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1235 = cs_196 ? vram16x16_2_io_portA_dout : _GEN_1231; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1236 = cs_196 | _GEN_1234; // @[MemMap.scala 108:16 110:18]
  wire  cs_197 = addr_230 >= 24'h981000 & addr_230 <= 24'h9817ff; // @[Util.scala 64:67]
  wire  _GEN_1237 = ~cpu_io_as ? 1'h0 : _GEN_1236; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1238 = cs_197 ? lineRam_2_io_portA_dout : _GEN_1235; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1239 = cs_197 | _GEN_1237; // @[MemMap.scala 108:16 110:18]
  wire  cs_198 = addr_230 >= 24'h981800 & addr_230 <= 24'h983fff; // @[Util.scala 64:67]
  wire  _GEN_1240 = ~cpu_io_as ? 1'h0 : _GEN_1239; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_34; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1242 = readStrobe ? tmp_34 : _GEN_1238; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1244 = cs_198 ? _GEN_1242 : _GEN_1238; // @[MemMap.scala 164:16]
  wire  _GEN_1246 = cs_198 | _GEN_1240; // @[MemMap.scala 164:16 170:18]
  wire  cs_199 = addr_230 >= 24'h984000 & addr_230 <= 24'h987fff; // @[Util.scala 64:67]
  wire  _GEN_1247 = ~cpu_io_as ? 1'h0 : _GEN_1246; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1248 = cs_199 ? vram8x8_2_io_portA_dout : _GEN_1244; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1249 = cs_199 | _GEN_1247; // @[MemMap.scala 108:16 110:18]
  wire  cs_200 = addr_230 >= 24'h988000 & addr_230 <= 24'h98ffff; // @[Util.scala 64:67]
  wire  _GEN_1250 = ~cpu_io_as ? 1'h0 : _GEN_1249; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_35; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1252 = readStrobe ? tmp_35 : _GEN_1248; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1254 = cs_200 ? _GEN_1252 : _GEN_1248; // @[MemMap.scala 164:16]
  wire  _GEN_1256 = cs_200 | _GEN_1250; // @[MemMap.scala 164:16 170:18]
  wire [23:0] offset_200 = addr_230 - 24'ha80000; // @[MemMap.scala 84:23]
  wire  cs_201 = addr_230 >= 24'ha80000 & addr_230 <= 24'ha80007; // @[Util.scala 64:67]
  wire  _GEN_1257 = ~cpu_io_as ? 1'h0 : _GEN_1256; // @[MemMap.scala 226:{19,30}]
  wire  dinReg_a_6 = offset_200 == 24'h0 & agalletIrq; // @[Main.scala 219:28]
  wire  _GEN_1258 = offset_200 == 24'h4 ? 1'h0 : _GEN_1111; // @[Main.scala 222:{26,37}]
  wire  _dinReg_T_38 = ~dinReg_a_6; // @[Main.scala 224:9]
  wire [2:0] _dinReg_T_41 = {_dinReg_T_38,1'h1,_dinReg_T_4}; // @[Cat.scala 33:92]
  wire  _GEN_1260 = cs_201 & readStrobe ? _GEN_1258 : _GEN_1111; // @[MemMap.scala 180:30]
  wire [15:0] _GEN_1262 = cs_201 & readStrobe ? {{13'd0}, _dinReg_T_41} : _GEN_1254; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_1263 = cs_201 & readStrobe | _GEN_1257; // @[MemMap.scala 180:30 182:18]
  wire  cs_202 = addr_230 >= 24'ha80000 & addr_230 <= 24'ha8000f; // @[Util.scala 64:67]
  wire  _GEN_1264 = ~cpu_io_as ? 1'h0 : _GEN_1263; // @[MemMap.scala 226:{19,30}]
  wire  mem_6_wr = cs_202 & writeStrobe; // @[MemMap.scala 150:20]
  wire  _GEN_1265 = cs_202 & _upperWriteStrobe_T_3 | _GEN_1264; // @[MemMap.scala 154:{27,38}]
  wire  cs_203 = addr_230 >= 24'ha80008 & addr_230 <= 24'ha80008; // @[Util.scala 64:67]
  wire  _GEN_1266 = ~cpu_io_as ? 1'h0 : _GEN_1265; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_1267 = cs_203 & writeStrobe | _GEN_1118; // @[MemMap.scala 192:31 Main.scala 258:68]
  wire  _GEN_1268 = cs_203 & writeStrobe | _GEN_1266; // @[MemMap.scala 192:31 194:18]
  wire  cs_204 = addr_230 >= 24'ha8000a & addr_230 <= 24'ha8007f; // @[Util.scala 64:67]
  wire  _GEN_1269 = ~cpu_io_as ? 1'h0 : _GEN_1268; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1270 = readStrobe ? 16'h0 : _GEN_1262; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1271 = cs_204 ? _GEN_1270 : _GEN_1262; // @[MemMap.scala 164:16]
  wire  _GEN_1272 = cs_204 | _GEN_1269; // @[MemMap.scala 164:16 170:18]
  wire  cs_205 = addr_230 >= 24'ha8006e & addr_230 <= 24'ha8006e; // @[Util.scala 64:67]
  wire  _GEN_1273 = ~cpu_io_as ? 1'h0 : _GEN_1272; // @[MemMap.scala 226:{19,30}]
  wire  _T_292 = cs_205 & writeStrobe; // @[MemMap.scala 192:15]
  wire  _GEN_1275 = cs_205 & writeStrobe | _GEN_1273; // @[MemMap.scala 192:31 194:18]
  wire  _GEN_1276 = ~cpu_io_as ? 1'h0 : _GEN_1275; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1277 = cs_77 ? layerRegs_0_io_mem_dout : _GEN_1271; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1278 = cs_77 | _GEN_1276; // @[MemMap.scala 108:16 110:18]
  wire  cs_207 = addr_230 >= 24'hb80000 & addr_230 <= 24'hb80005; // @[Util.scala 64:67]
  wire  _GEN_1279 = ~cpu_io_as ? 1'h0 : _GEN_1278; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1280 = cs_207 ? layerRegs_1_io_mem_dout : _GEN_1277; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1281 = cs_207 | _GEN_1279; // @[MemMap.scala 108:16 110:18]
  wire  cs_208 = addr_230 >= 24'hc00000 & addr_230 <= 24'hc00005; // @[Util.scala 64:67]
  wire  _GEN_1282 = ~cpu_io_as ? 1'h0 : _GEN_1281; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1283 = cs_208 ? layerRegs_2_io_mem_dout : _GEN_1280; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1284 = cs_208 | _GEN_1282; // @[MemMap.scala 108:16 110:18]
  wire  cs_209 = addr_230 >= 24'hc80000 & addr_230 <= 24'hc80000; // @[Util.scala 64:67]
  wire  _GEN_1285 = ~cpu_io_as ? 1'h0 : _GEN_1284; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1286 = cs_209 & readStrobe ? input0 : _GEN_1283; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_1287 = cs_209 & readStrobe | _GEN_1285; // @[MemMap.scala 180:30 182:18]
  wire  cs_210 = addr_230 >= 24'hc80002 & addr_230 <= 24'hc80002; // @[Util.scala 64:67]
  wire  _GEN_1288 = ~cpu_io_as ? 1'h0 : _GEN_1287; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1289 = cs_210 & readStrobe ? input1 : _GEN_1286; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_1290 = cs_210 & readStrobe | _GEN_1288; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_1291 = ~cpu_io_as ? 1'h0 : _GEN_1290; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_1292 = cs_211 & _upperWriteStrobe_T_3 | _GEN_1291; // @[MemMap.scala 154:{27,38}]
  wire  _GEN_1293 = ~cpu_io_as ? 1'h0 : _GEN_1292; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1294 = readStrobe ? 16'h0 : _GEN_1289; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1295 = cs_80 ? _GEN_1294 : _GEN_1289; // @[MemMap.scala 164:16]
  wire  _GEN_1296 = cs_80 | _GEN_1293; // @[MemMap.scala 164:16 170:18]
  wire  cs_213 = addr_230 >= 24'hf00000 & addr_230 <= 24'hf0ffff; // @[Util.scala 64:67]
  wire  _GEN_1297 = ~cpu_io_as ? 1'h0 : _GEN_1296; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1298 = cs_213 ? spriteRam_io_portA_dout : _GEN_1295; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1299 = cs_213 | _GEN_1297; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1300 = io_gameIndex == 4'h7 ? _GEN_1299 : _GEN_1100; // @[Main.scala 393:42]
  wire  _GEN_1303 = io_gameIndex == 4'h7 ? cs_2 & readStrobe : _GEN_1103; // @[Main.scala 393:42 MemMap.scala 128:14]
  wire [23:0] _GEN_1304 = io_gameIndex == 4'h7 ? addr_230 : _GEN_1104; // @[Main.scala 393:42 MemMap.scala 129:16]
  wire [15:0] _GEN_1305 = io_gameIndex == 4'h7 ? _GEN_1298 : _GEN_1105; // @[Main.scala 393:42]
  wire  _GEN_1306 = io_gameIndex == 4'h7 ? cs_183 & readStrobe : _GEN_1106; // @[Main.scala 393:42 MemMap.scala 103:14]
  wire  _GEN_1307 = io_gameIndex == 4'h7 ? cs_183 & writeStrobe : _GEN_1107; // @[Main.scala 393:42 MemMap.scala 104:14]
  wire [22:0] _GEN_1308 = io_gameIndex == 4'h7 ? cpu_io_addr : _GEN_1108; // @[Main.scala 393:42 MemMap.scala 105:16]
  wire [1:0] _GEN_1309 = io_gameIndex == 4'h7 ? _mainRam_io_mask_T : _GEN_1109; // @[Main.scala 393:42 MemMap.scala 106:16]
  wire [15:0] _GEN_1310 = io_gameIndex == 4'h7 ? cpu_io_dout : _GEN_1110; // @[Main.scala 393:42 MemMap.scala 107:15]
  wire  _GEN_1311 = io_gameIndex == 4'h7 ? cs_184 & readStrobe : _GEN_1168; // @[Main.scala 393:42 MemMap.scala 103:14]
  wire  _GEN_1312 = io_gameIndex == 4'h7 ? cs_184 & writeStrobe : _GEN_1169; // @[Main.scala 393:42 MemMap.scala 104:14]
  wire [22:0] _GEN_1313 = io_gameIndex == 4'h7 ? {{12'd0}, cpu_io_addr[10:0]} : _GEN_1170; // @[Main.scala 393:42 MemMap.scala 105:16]
  wire  _GEN_1315 = io_gameIndex == 4'h7 ? cs_186 & readStrobe : _GEN_1122; // @[Main.scala 393:42 MemMap.scala 103:14]
  wire  _GEN_1316 = io_gameIndex == 4'h7 ? cs_186 & writeStrobe : _GEN_1123; // @[Main.scala 393:42 MemMap.scala 104:14]
  wire  _GEN_1318 = io_gameIndex == 4'h7 ? cs_187 & readStrobe : _GEN_1125; // @[Main.scala 393:42 MemMap.scala 103:14]
  wire  _GEN_1319 = io_gameIndex == 4'h7 ? cs_187 & writeStrobe : _GEN_1126; // @[Main.scala 393:42 MemMap.scala 104:14]
  wire  _GEN_1321 = io_gameIndex == 4'h7 ? cs_189 & readStrobe : _GEN_1128; // @[Main.scala 393:42 MemMap.scala 103:14]
  wire  _GEN_1322 = io_gameIndex == 4'h7 ? cs_189 & writeStrobe : _GEN_1129; // @[Main.scala 393:42 MemMap.scala 104:14]
  wire [22:0] _GEN_1335 = io_gameIndex == 4'h7 ? cpu_io_addr : _GEN_1142; // @[Main.scala 393:42 MemMap.scala 105:16]
  wire [22:0] _GEN_1343 = io_gameIndex == 4'h7 ? cpu_io_addr : _GEN_1150; // @[Main.scala 393:42 MemMap.scala 105:16]
  wire  _GEN_1346 = io_gameIndex == 4'h7 ? _GEN_1260 : _GEN_1111; // @[Main.scala 393:42]
  wire  _GEN_1349 = io_gameIndex == 4'h7 ? mem_6_wr : _GEN_1114; // @[Main.scala 393:42 MemIO.scala 305:8]
  wire [2:0] _GEN_1350 = io_gameIndex == 4'h7 ? mem_addr : _GEN_1115; // @[Main.scala 393:42 MemIO.scala 306:10]
  wire [15:0] _GEN_1352 = io_gameIndex == 4'h7 ? _GEN_193 : _GEN_1117; // @[Main.scala 393:42 MemIO.scala 308:9]
  wire  _GEN_1353 = io_gameIndex == 4'h7 ? _GEN_1267 : _GEN_1118; // @[Main.scala 393:42]
  wire  _GEN_1356 = io_gameIndex == 4'h7 ? cs_77 & writeStrobe : _GEN_1159; // @[Main.scala 393:42 MemMap.scala 104:14]
  wire [22:0] _GEN_1363 = io_gameIndex == 4'h7 ? cpu_io_addr : _GEN_1155; // @[Main.scala 393:42 MemMap.scala 105:16]
  wire  _GEN_1369 = io_gameIndex == 4'h7 ? cs_213 & readStrobe : _GEN_1119; // @[Main.scala 393:42 MemMap.scala 103:14]
  wire  _GEN_1370 = io_gameIndex == 4'h7 ? cs_213 & writeStrobe : _GEN_1120; // @[Main.scala 393:42 MemMap.scala 104:14]
  wire  _GEN_1372 = ~cpu_io_as ? 1'h0 : _GEN_1300; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1373 = cs_2 & cpu_io_rw & io_progRom_valid ? io_progRom_dout : _GEN_1305; // @[MemMap.scala 130:39 131:16]
  wire  _GEN_1374 = cs_2 & cpu_io_rw & io_progRom_valid | _GEN_1372; // @[MemMap.scala 130:39 132:18]
  wire  _GEN_1375 = ~cpu_io_as ? 1'h0 : _GEN_1374; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1376 = cs_3 ? mainRam_io_dout : _GEN_1373; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1377 = cs_3 | _GEN_1375; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1378 = ~cpu_io_as ? 1'h0 : _GEN_1377; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1379 = cs_4 ? io_soundCtrl_ymz_dout : _GEN_1376; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1380 = cs_4 | _GEN_1378; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1381 = ~cpu_io_as ? 1'h0 : _GEN_1380; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1382 = cs_5 ? spriteRam_io_portA_dout : _GEN_1379; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1383 = cs_5 | _GEN_1381; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1384 = ~cpu_io_as ? 1'h0 : _GEN_1383; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1385 = cs_6 ? vram16x16_0_io_portA_dout : _GEN_1382; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1386 = cs_6 | _GEN_1384; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1387 = ~cpu_io_as ? 1'h0 : _GEN_1386; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1388 = cs_7 ? lineRam_0_io_portA_dout : _GEN_1385; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1389 = cs_7 | _GEN_1387; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1390 = ~cpu_io_as ? 1'h0 : _GEN_1389; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_36; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1392 = readStrobe ? tmp_36 : _GEN_1388; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1394 = cs_8 ? _GEN_1392 : _GEN_1388; // @[MemMap.scala 164:16]
  wire  _GEN_1396 = cs_8 | _GEN_1390; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_1397 = ~cpu_io_as ? 1'h0 : _GEN_1396; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1398 = cs_9 ? vram8x8_0_io_portA_dout : _GEN_1394; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1399 = cs_9 | _GEN_1397; // @[MemMap.scala 108:16 110:18]
  wire  _GEN_1400 = ~cpu_io_as ? 1'h0 : _GEN_1399; // @[MemMap.scala 226:{19,30}]
  reg [15:0] tmp_37; // @[MemMap.scala 206:20]
  wire [15:0] _GEN_1402 = readStrobe ? tmp_37 : _GEN_1398; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1404 = cs_10 ? _GEN_1402 : _GEN_1398; // @[MemMap.scala 164:16]
  wire  _GEN_1406 = cs_10 | _GEN_1400; // @[MemMap.scala 164:16 170:18]
  wire  cs_223 = addr_230 >= 24'h600000 & addr_230 <= 24'h600007; // @[Util.scala 64:67]
  wire  _GEN_1407 = ~cpu_io_as ? 1'h0 : _GEN_1406; // @[MemMap.scala 226:{19,30}]
  wire  dinReg_a_7 = offset_10 == 24'h0 & agalletIrq; // @[Main.scala 219:28]
  wire  _dinReg_T_44 = ~dinReg_a_7; // @[Main.scala 224:9]
  wire [2:0] _dinReg_T_47 = {_dinReg_T_44,1'h1,_dinReg_T_4}; // @[Cat.scala 33:92]
  wire [15:0] _GEN_1412 = cs_223 & readStrobe ? {{13'd0}, _dinReg_T_47} : _GEN_1404; // @[MemMap.scala 180:30 181:16]
  wire  _GEN_1413 = cs_223 & readStrobe | _GEN_1407; // @[MemMap.scala 180:30 182:18]
  wire  cs_224 = addr_230 >= 24'h600000 & addr_230 <= 24'h60000f; // @[Util.scala 64:67]
  wire  _GEN_1414 = ~cpu_io_as ? 1'h0 : _GEN_1413; // @[MemMap.scala 226:{19,30}]
  wire  mem_7_wr = cs_224 & writeStrobe; // @[MemMap.scala 150:20]
  wire  _GEN_1415 = cs_224 & _upperWriteStrobe_T_3 | _GEN_1414; // @[MemMap.scala 154:{27,38}]
  wire  cs_225 = addr_230 >= 24'h600008 & addr_230 <= 24'h600008; // @[Util.scala 64:67]
  wire  _GEN_1416 = ~cpu_io_as ? 1'h0 : _GEN_1415; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_1417 = cs_225 & writeStrobe | _GEN_1353; // @[MemMap.scala 192:31 Main.scala 258:68]
  wire  _GEN_1418 = cs_225 & writeStrobe | _GEN_1416; // @[MemMap.scala 192:31 194:18]
  wire  cs_226 = addr_230 >= 24'h60000a & addr_230 <= 24'h60007f; // @[Util.scala 64:67]
  wire  _GEN_1419 = ~cpu_io_as ? 1'h0 : _GEN_1418; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1420 = readStrobe ? 16'h0 : _GEN_1412; // @[MemMap.scala 165:26 166:18]
  wire [15:0] _GEN_1421 = cs_226 ? _GEN_1420 : _GEN_1412; // @[MemMap.scala 164:16]
  wire  _GEN_1422 = cs_226 | _GEN_1419; // @[MemMap.scala 164:16 170:18]
  wire  _GEN_1423 = ~cpu_io_as ? 1'h0 : _GEN_1422; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1424 = cs_42 ? layerRegs_0_io_mem_dout : _GEN_1421; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1425 = cs_42 | _GEN_1423; // @[MemMap.scala 108:16 110:18]
  wire  cs_228 = addr_230 >= 24'h800000 & addr_230 <= 24'h80ffff; // @[Util.scala 64:67]
  wire  _GEN_1426 = ~cpu_io_as ? 1'h0 : _GEN_1425; // @[MemMap.scala 226:{19,30}]
  wire [15:0] _GEN_1427 = cs_228 ? paletteRam_io_portA_dout : _GEN_1424; // @[MemMap.scala 108:16 109:16]
  wire  _GEN_1428 = cs_228 | _GEN_1426; // @[MemMap.scala 108:16 110:18]
  wire  cs_229 = addr_230 >= 24'h900000 & addr_230 <= 24'h900000; // @[Util.scala 64:67]
  wire  _GEN_1429 = ~cpu_io_as ? 1'h0 : _GEN_1428; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_1431 = cs_229 & readStrobe | _GEN_1429; // @[MemMap.scala 180:30 182:18]
  wire  cs_230 = addr_230 >= 24'h900002 & addr_230 <= 24'h900002; // @[Util.scala 64:67]
  wire  _GEN_1432 = ~cpu_io_as ? 1'h0 : _GEN_1431; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_1434 = cs_230 & readStrobe | _GEN_1432; // @[MemMap.scala 180:30 182:18]
  wire  _GEN_1435 = ~cpu_io_as ? 1'h0 : _GEN_1434; // @[MemMap.scala 226:{19,30}]
  wire  _GEN_1436 = cs_231 & _upperWriteStrobe_T_3 | _GEN_1435; // @[MemMap.scala 154:{27,38}]
  wire [23:0] _GEN_1441 = io_gameIndex == 4'h4 ? addr_230 : _GEN_1304; // @[Main.scala 414:40 MemMap.scala 129:16]
  wire [22:0] _GEN_1445 = io_gameIndex == 4'h4 ? cpu_io_addr : _GEN_1308; // @[Main.scala 414:40 MemMap.scala 105:16]
  wire [22:0] _GEN_1478 = io_gameIndex == 4'h4 ? cpu_io_addr : _GEN_1313; // @[Main.scala 414:40 MemMap.scala 105:16]
  CPU cpu ( // @[Main.scala 91:19]
    .clock(cpu_clock),
    .reset(cpu_reset),
    .io_halt(cpu_io_halt),
    .io_as(cpu_io_as),
    .io_rw(cpu_io_rw),
    .io_uds(cpu_io_uds),
    .io_lds(cpu_io_lds),
    .io_dtack(cpu_io_dtack),
    .io_vpa(cpu_io_vpa),
    .io_ipl(cpu_io_ipl),
    .io_fc(cpu_io_fc),
    .io_addr(cpu_io_addr),
    .io_din(cpu_io_din),
    .io_dout(cpu_io_dout)
  );
  EEPROM eeprom ( // @[Main.scala 109:22]
    .clock(eeprom_clock),
    .reset(eeprom_reset),
    .io_mem_rd(eeprom_io_mem_rd),
    .io_mem_wr(eeprom_io_mem_wr),
    .io_mem_addr(eeprom_io_mem_addr),
    .io_mem_din(eeprom_io_mem_din),
    .io_mem_dout(eeprom_io_mem_dout),
    .io_mem_wait_n(eeprom_io_mem_wait_n),
    .io_mem_valid(eeprom_io_mem_valid),
    .io_serial_cs(eeprom_io_serial_cs),
    .io_serial_sck(eeprom_io_serial_sck),
    .io_serial_sdi(eeprom_io_serial_sdi),
    .io_serial_sdo(eeprom_io_serial_sdo)
  );
  SinglePortRam mainRam ( // @[Main.scala 120:23]
    .clock(mainRam_clock),
    .io_rd(mainRam_io_rd),
    .io_wr(mainRam_io_wr),
    .io_addr(mainRam_io_addr),
    .io_mask(mainRam_io_mask),
    .io_din(mainRam_io_din),
    .io_dout(mainRam_io_dout)
  );
  TrueDualPortRam spriteRam ( // @[Main.scala 128:25]
    .clock(spriteRam_clock),
    .io_clockB(spriteRam_io_clockB),
    .io_portA_rd(spriteRam_io_portA_rd),
    .io_portA_wr(spriteRam_io_portA_wr),
    .io_portA_addr(spriteRam_io_portA_addr),
    .io_portA_mask(spriteRam_io_portA_mask),
    .io_portA_din(spriteRam_io_portA_din),
    .io_portA_dout(spriteRam_io_portA_dout),
    .io_portB_rd(spriteRam_io_portB_rd),
    .io_portB_addr(spriteRam_io_portB_addr),
    .io_portB_dout(spriteRam_io_portB_dout)
  );
  TrueDualPortRam_1 vram8x8_0 ( // @[Main.scala 141:21]
    .clock(vram8x8_0_clock),
    .io_clockB(vram8x8_0_io_clockB),
    .io_portA_rd(vram8x8_0_io_portA_rd),
    .io_portA_wr(vram8x8_0_io_portA_wr),
    .io_portA_addr(vram8x8_0_io_portA_addr),
    .io_portA_mask(vram8x8_0_io_portA_mask),
    .io_portA_din(vram8x8_0_io_portA_din),
    .io_portA_dout(vram8x8_0_io_portA_dout),
    .io_portB_addr(vram8x8_0_io_portB_addr),
    .io_portB_dout(vram8x8_0_io_portB_dout)
  );
  TrueDualPortRam_1 vram8x8_1 ( // @[Main.scala 141:21]
    .clock(vram8x8_1_clock),
    .io_clockB(vram8x8_1_io_clockB),
    .io_portA_rd(vram8x8_1_io_portA_rd),
    .io_portA_wr(vram8x8_1_io_portA_wr),
    .io_portA_addr(vram8x8_1_io_portA_addr),
    .io_portA_mask(vram8x8_1_io_portA_mask),
    .io_portA_din(vram8x8_1_io_portA_din),
    .io_portA_dout(vram8x8_1_io_portA_dout),
    .io_portB_addr(vram8x8_1_io_portB_addr),
    .io_portB_dout(vram8x8_1_io_portB_dout)
  );
  TrueDualPortRam_1 vram8x8_2 ( // @[Main.scala 141:21]
    .clock(vram8x8_2_clock),
    .io_clockB(vram8x8_2_io_clockB),
    .io_portA_rd(vram8x8_2_io_portA_rd),
    .io_portA_wr(vram8x8_2_io_portA_wr),
    .io_portA_addr(vram8x8_2_io_portA_addr),
    .io_portA_mask(vram8x8_2_io_portA_mask),
    .io_portA_din(vram8x8_2_io_portA_din),
    .io_portA_dout(vram8x8_2_io_portA_dout),
    .io_portB_addr(vram8x8_2_io_portB_addr),
    .io_portB_dout(vram8x8_2_io_portB_dout)
  );
  TrueDualPortRam_4 vram16x16_0 ( // @[Main.scala 156:21]
    .clock(vram16x16_0_clock),
    .io_clockB(vram16x16_0_io_clockB),
    .io_portA_rd(vram16x16_0_io_portA_rd),
    .io_portA_wr(vram16x16_0_io_portA_wr),
    .io_portA_addr(vram16x16_0_io_portA_addr),
    .io_portA_mask(vram16x16_0_io_portA_mask),
    .io_portA_din(vram16x16_0_io_portA_din),
    .io_portA_dout(vram16x16_0_io_portA_dout),
    .io_portB_addr(vram16x16_0_io_portB_addr),
    .io_portB_dout(vram16x16_0_io_portB_dout)
  );
  TrueDualPortRam_4 vram16x16_1 ( // @[Main.scala 156:21]
    .clock(vram16x16_1_clock),
    .io_clockB(vram16x16_1_io_clockB),
    .io_portA_rd(vram16x16_1_io_portA_rd),
    .io_portA_wr(vram16x16_1_io_portA_wr),
    .io_portA_addr(vram16x16_1_io_portA_addr),
    .io_portA_mask(vram16x16_1_io_portA_mask),
    .io_portA_din(vram16x16_1_io_portA_din),
    .io_portA_dout(vram16x16_1_io_portA_dout),
    .io_portB_addr(vram16x16_1_io_portB_addr),
    .io_portB_dout(vram16x16_1_io_portB_dout)
  );
  TrueDualPortRam_4 vram16x16_2 ( // @[Main.scala 156:21]
    .clock(vram16x16_2_clock),
    .io_clockB(vram16x16_2_io_clockB),
    .io_portA_rd(vram16x16_2_io_portA_rd),
    .io_portA_wr(vram16x16_2_io_portA_wr),
    .io_portA_addr(vram16x16_2_io_portA_addr),
    .io_portA_mask(vram16x16_2_io_portA_mask),
    .io_portA_din(vram16x16_2_io_portA_din),
    .io_portA_dout(vram16x16_2_io_portA_dout),
    .io_portB_addr(vram16x16_2_io_portB_addr),
    .io_portB_dout(vram16x16_2_io_portB_dout)
  );
  TrueDualPortRam_7 lineRam_0 ( // @[Main.scala 171:21]
    .clock(lineRam_0_clock),
    .io_clockB(lineRam_0_io_clockB),
    .io_portA_rd(lineRam_0_io_portA_rd),
    .io_portA_wr(lineRam_0_io_portA_wr),
    .io_portA_addr(lineRam_0_io_portA_addr),
    .io_portA_mask(lineRam_0_io_portA_mask),
    .io_portA_din(lineRam_0_io_portA_din),
    .io_portA_dout(lineRam_0_io_portA_dout),
    .io_portB_addr(lineRam_0_io_portB_addr),
    .io_portB_dout(lineRam_0_io_portB_dout)
  );
  TrueDualPortRam_7 lineRam_1 ( // @[Main.scala 171:21]
    .clock(lineRam_1_clock),
    .io_clockB(lineRam_1_io_clockB),
    .io_portA_rd(lineRam_1_io_portA_rd),
    .io_portA_wr(lineRam_1_io_portA_wr),
    .io_portA_addr(lineRam_1_io_portA_addr),
    .io_portA_mask(lineRam_1_io_portA_mask),
    .io_portA_din(lineRam_1_io_portA_din),
    .io_portA_dout(lineRam_1_io_portA_dout),
    .io_portB_addr(lineRam_1_io_portB_addr),
    .io_portB_dout(lineRam_1_io_portB_dout)
  );
  TrueDualPortRam_7 lineRam_2 ( // @[Main.scala 171:21]
    .clock(lineRam_2_clock),
    .io_clockB(lineRam_2_io_clockB),
    .io_portA_rd(lineRam_2_io_portA_rd),
    .io_portA_wr(lineRam_2_io_portA_wr),
    .io_portA_addr(lineRam_2_io_portA_addr),
    .io_portA_mask(lineRam_2_io_portA_mask),
    .io_portA_din(lineRam_2_io_portA_din),
    .io_portA_dout(lineRam_2_io_portA_dout),
    .io_portB_addr(lineRam_2_io_portB_addr),
    .io_portB_dout(lineRam_2_io_portB_dout)
  );
  TrueDualPortRam_10 paletteRam ( // @[Main.scala 185:26]
    .clock(paletteRam_clock),
    .io_clockB(paletteRam_io_clockB),
    .io_portA_rd(paletteRam_io_portA_rd),
    .io_portA_wr(paletteRam_io_portA_wr),
    .io_portA_addr(paletteRam_io_portA_addr),
    .io_portA_mask(paletteRam_io_portA_mask),
    .io_portA_din(paletteRam_io_portA_din),
    .io_portA_dout(paletteRam_io_portA_dout),
    .io_portB_addr(paletteRam_io_portB_addr),
    .io_portB_dout(paletteRam_io_portB_dout)
  );
  RegisterFile_2 layerRegs_0 ( // @[Main.scala 198:22]
    .clock(layerRegs_0_clock),
    .io_mem_wr(layerRegs_0_io_mem_wr),
    .io_mem_addr(layerRegs_0_io_mem_addr),
    .io_mem_mask(layerRegs_0_io_mem_mask),
    .io_mem_din(layerRegs_0_io_mem_din),
    .io_mem_dout(layerRegs_0_io_mem_dout),
    .io_regs_0(layerRegs_0_io_regs_0),
    .io_regs_1(layerRegs_0_io_regs_1),
    .io_regs_2(layerRegs_0_io_regs_2)
  );
  RegisterFile_2 layerRegs_1 ( // @[Main.scala 198:22]
    .clock(layerRegs_1_clock),
    .io_mem_wr(layerRegs_1_io_mem_wr),
    .io_mem_addr(layerRegs_1_io_mem_addr),
    .io_mem_mask(layerRegs_1_io_mem_mask),
    .io_mem_din(layerRegs_1_io_mem_din),
    .io_mem_dout(layerRegs_1_io_mem_dout),
    .io_regs_0(layerRegs_1_io_regs_0),
    .io_regs_1(layerRegs_1_io_regs_1),
    .io_regs_2(layerRegs_1_io_regs_2)
  );
  RegisterFile_2 layerRegs_2 ( // @[Main.scala 198:22]
    .clock(layerRegs_2_clock),
    .io_mem_wr(layerRegs_2_io_mem_wr),
    .io_mem_addr(layerRegs_2_io_mem_addr),
    .io_mem_mask(layerRegs_2_io_mem_mask),
    .io_mem_din(layerRegs_2_io_mem_din),
    .io_mem_dout(layerRegs_2_io_mem_dout),
    .io_regs_0(layerRegs_2_io_regs_0),
    .io_regs_1(layerRegs_2_io_regs_1),
    .io_regs_2(layerRegs_2_io_regs_2)
  );
  RegisterFile_5 spriteRegs ( // @[Main.scala 205:26]
    .clock(spriteRegs_clock),
    .io_mem_wr(spriteRegs_io_mem_wr),
    .io_mem_addr(spriteRegs_io_mem_addr),
    .io_mem_mask(spriteRegs_io_mem_mask),
    .io_mem_din(spriteRegs_io_mem_din),
    .io_regs_0(spriteRegs_io_regs_0),
    .io_regs_1(spriteRegs_io_regs_1),
    .io_regs_4(spriteRegs_io_regs_4),
    .io_regs_5(spriteRegs_io_regs_5)
  );
  assign io_gpuMem_layer_0_regs_tileSize = io_gpuMem_layer_0_regs_r_1_tileSize; // @[Main.scala 200:29]
  assign io_gpuMem_layer_0_regs_enable = io_gpuMem_layer_0_regs_r_1_enable; // @[Main.scala 200:29]
  assign io_gpuMem_layer_0_regs_flipX = io_gpuMem_layer_0_regs_r_1_flipX; // @[Main.scala 200:29]
  assign io_gpuMem_layer_0_regs_flipY = io_gpuMem_layer_0_regs_r_1_flipY; // @[Main.scala 200:29]
  assign io_gpuMem_layer_0_regs_rowScrollEnable = io_gpuMem_layer_0_regs_r_1_rowScrollEnable; // @[Main.scala 200:29]
  assign io_gpuMem_layer_0_regs_rowSelectEnable = io_gpuMem_layer_0_regs_r_1_rowSelectEnable; // @[Main.scala 200:29]
  assign io_gpuMem_layer_0_regs_scroll_x = io_gpuMem_layer_0_regs_r_1_scroll_x; // @[Main.scala 200:29]
  assign io_gpuMem_layer_0_regs_scroll_y = io_gpuMem_layer_0_regs_r_1_scroll_y; // @[Main.scala 200:29]
  assign io_gpuMem_layer_0_vram8x8_dout = vram8x8_0_io_portB_dout; // @[Main.scala 150:18]
  assign io_gpuMem_layer_0_vram16x16_dout = vram16x16_0_io_portB_dout; // @[Main.scala 165:18]
  assign io_gpuMem_layer_0_lineRam_dout = lineRam_0_io_portB_dout; // @[Main.scala 180:18]
  assign io_gpuMem_layer_1_regs_tileSize = io_gpuMem_layer_1_regs_r_1_tileSize; // @[Main.scala 200:29]
  assign io_gpuMem_layer_1_regs_enable = io_gpuMem_layer_1_regs_r_1_enable; // @[Main.scala 200:29]
  assign io_gpuMem_layer_1_regs_flipX = io_gpuMem_layer_1_regs_r_1_flipX; // @[Main.scala 200:29]
  assign io_gpuMem_layer_1_regs_flipY = io_gpuMem_layer_1_regs_r_1_flipY; // @[Main.scala 200:29]
  assign io_gpuMem_layer_1_regs_rowScrollEnable = io_gpuMem_layer_1_regs_r_1_rowScrollEnable; // @[Main.scala 200:29]
  assign io_gpuMem_layer_1_regs_rowSelectEnable = io_gpuMem_layer_1_regs_r_1_rowSelectEnable; // @[Main.scala 200:29]
  assign io_gpuMem_layer_1_regs_scroll_x = io_gpuMem_layer_1_regs_r_1_scroll_x; // @[Main.scala 200:29]
  assign io_gpuMem_layer_1_regs_scroll_y = io_gpuMem_layer_1_regs_r_1_scroll_y; // @[Main.scala 200:29]
  assign io_gpuMem_layer_1_vram8x8_dout = vram8x8_1_io_portB_dout; // @[Main.scala 150:18]
  assign io_gpuMem_layer_1_vram16x16_dout = vram16x16_1_io_portB_dout; // @[Main.scala 165:18]
  assign io_gpuMem_layer_1_lineRam_dout = lineRam_1_io_portB_dout; // @[Main.scala 180:18]
  assign io_gpuMem_layer_2_regs_tileSize = io_gpuMem_layer_2_regs_r_1_tileSize; // @[Main.scala 200:29]
  assign io_gpuMem_layer_2_regs_enable = io_gpuMem_layer_2_regs_r_1_enable; // @[Main.scala 200:29]
  assign io_gpuMem_layer_2_regs_flipX = io_gpuMem_layer_2_regs_r_1_flipX; // @[Main.scala 200:29]
  assign io_gpuMem_layer_2_regs_flipY = io_gpuMem_layer_2_regs_r_1_flipY; // @[Main.scala 200:29]
  assign io_gpuMem_layer_2_regs_rowScrollEnable = io_gpuMem_layer_2_regs_r_1_rowScrollEnable; // @[Main.scala 200:29]
  assign io_gpuMem_layer_2_regs_rowSelectEnable = io_gpuMem_layer_2_regs_r_1_rowSelectEnable; // @[Main.scala 200:29]
  assign io_gpuMem_layer_2_regs_scroll_x = io_gpuMem_layer_2_regs_r_1_scroll_x; // @[Main.scala 200:29]
  assign io_gpuMem_layer_2_regs_scroll_y = io_gpuMem_layer_2_regs_r_1_scroll_y; // @[Main.scala 200:29]
  assign io_gpuMem_layer_2_vram8x8_dout = vram8x8_2_io_portB_dout; // @[Main.scala 150:18]
  assign io_gpuMem_layer_2_vram16x16_dout = vram16x16_2_io_portB_dout; // @[Main.scala 165:18]
  assign io_gpuMem_layer_2_lineRam_dout = lineRam_2_io_portB_dout; // @[Main.scala 180:18]
  assign io_gpuMem_sprite_regs_offset_x = spriteRegs_io_regs_0[8:0]; // @[SpriteRegs.scala 78:33]
  assign io_gpuMem_sprite_regs_offset_y = spriteRegs_io_regs_1[8:0]; // @[SpriteRegs.scala 78:48]
  assign io_gpuMem_sprite_regs_bank = spriteRegs_io_regs_4[1:0]; // @[SpriteRegs.scala 79:25]
  assign io_gpuMem_sprite_regs_fixed = |spriteRegs_io_regs_5[13:12]; // @[SpriteRegs.scala 80:35]
  assign io_gpuMem_sprite_regs_hFlip = spriteRegs_io_regs_0[15]; // @[SpriteRegs.scala 76:26]
  assign io_gpuMem_sprite_vram_dout = spriteRam_io_portB_dout; // @[Main.scala 137:22]
  assign io_gpuMem_paletteRam_dout = paletteRam_io_portB_dout; // @[Main.scala 194:23]
  assign io_soundCtrl_oki_0_wr = io_gameIndex == 4'h2 & (cs_49 & writeStrobe); // @[Main.scala 285:42 MemMap.scala 104:14 MemIO.scala 318:8]
  assign io_soundCtrl_oki_0_din = cpu_io_dout; // @[Main.scala 285:42 MemMap.scala 107:15]
  assign io_soundCtrl_oki_1_wr = io_gameIndex == 4'h2 & (cs_50 & writeStrobe); // @[Main.scala 285:42 MemMap.scala 104:14 MemIO.scala 318:8]
  assign io_soundCtrl_oki_1_din = cpu_io_dout; // @[Main.scala 285:42 MemMap.scala 107:15]
  assign io_soundCtrl_nmk_wr = io_gameIndex == 4'h2 & (cs_51 & writeStrobe); // @[Main.scala 285:42 MemMap.scala 150:14 MemIO.scala 207:8]
  assign io_soundCtrl_nmk_addr = cpu_io_addr; // @[Main.scala 285:42 MemMap.scala 105:16]
  assign io_soundCtrl_nmk_din = cpu_io_dout; // @[Main.scala 285:42 MemMap.scala 107:15]
  assign io_soundCtrl_ymz_rd = io_gameIndex == 4'h4 ? cs_4 & readStrobe : _GEN_1153; // @[Main.scala 414:40 MemMap.scala 103:14]
  assign io_soundCtrl_ymz_wr = io_gameIndex == 4'h4 ? cs_4 & writeStrobe : _GEN_1154; // @[Main.scala 414:40 MemMap.scala 104:14]
  assign io_soundCtrl_ymz_addr = io_gameIndex == 4'h4 ? cpu_io_addr : _GEN_1155; // @[Main.scala 414:40 MemMap.scala 105:16]
  assign io_soundCtrl_ymz_din = io_gameIndex == 4'h4 ? cpu_io_dout : _GEN_1152; // @[Main.scala 414:40 MemMap.scala 107:15]
  assign io_soundCtrl_req = io_gameIndex == 4'h7 & _T_292; // @[Main.scala 104:20 393:42]
  assign io_soundCtrl_data = cpu_io_dout; // @[Main.scala 105:21]
  assign io_progRom_rd = io_gameIndex == 4'h4 ? cs_2 & readStrobe : _GEN_1303; // @[Main.scala 414:40 MemMap.scala 128:14]
  assign io_progRom_addr = _GEN_1441[19:0];
  assign io_eeprom_rd = eeprom_io_mem_rd; // @[Main.scala 110:17]
  assign io_eeprom_wr = eeprom_io_mem_wr; // @[Main.scala 110:17]
  assign io_eeprom_addr = eeprom_io_mem_addr; // @[Main.scala 110:17]
  assign io_eeprom_din = eeprom_io_mem_din; // @[Main.scala 110:17]
  assign io_spriteFrameBufferSwap = io_gameIndex == 4'h4 ? _GEN_1417 : _GEN_1353; // @[Main.scala 414:40]
  assign cpu_clock = clock;
  assign cpu_reset = reset;
  assign cpu_io_halt = pauseReg; // @[Main.scala 93:15]
  assign cpu_io_dtack = dtackReg; // @[Main.scala 414:40 MemMap.scala 230:15]
  assign cpu_io_vpa = cpu_io_as & cpu_io_fc == 3'h7; // @[Main.scala 95:27]
  assign cpu_io_ipl = {{2'd0}, _cpu_io_ipl_T}; // @[Main.scala 96:14]
  assign cpu_io_din = dinReg; // @[Main.scala 414:40 MemMap.scala 229:13]
  assign eeprom_clock = clock;
  assign eeprom_reset = reset;
  assign eeprom_io_mem_dout = io_eeprom_dout; // @[Main.scala 110:17]
  assign eeprom_io_mem_wait_n = io_eeprom_wait_n; // @[Main.scala 110:17]
  assign eeprom_io_mem_valid = io_eeprom_valid; // @[Main.scala 110:17]
  assign eeprom_io_serial_cs = eeprom_io_serial_cs_r; // @[Main.scala 114:23]
  assign eeprom_io_serial_sck = eeprom_io_serial_sck_r; // @[Main.scala 115:24]
  assign eeprom_io_serial_sdi = eeprom_io_serial_sdi_r; // @[Main.scala 116:24]
  assign mainRam_clock = clock;
  assign mainRam_io_rd = io_gameIndex == 4'h4 ? cs_3 & readStrobe : _GEN_1306; // @[Main.scala 414:40 MemMap.scala 103:14]
  assign mainRam_io_wr = io_gameIndex == 4'h4 ? cs_3 & writeStrobe : _GEN_1307; // @[Main.scala 414:40 MemMap.scala 104:14]
  assign mainRam_io_addr = _GEN_1445[14:0];
  assign mainRam_io_mask = io_gameIndex == 4'h4 ? _mainRam_io_mask_T : _GEN_1309; // @[Main.scala 414:40 MemMap.scala 106:16]
  assign mainRam_io_din = io_gameIndex == 4'h4 ? cpu_io_dout : _GEN_1310; // @[Main.scala 414:40 MemMap.scala 107:15]
  assign spriteRam_clock = clock;
  assign spriteRam_io_clockB = io_spriteClock; // @[Main.scala 135:23]
  assign spriteRam_io_portA_rd = io_gameIndex == 4'h4 ? cs_5 & readStrobe : _GEN_1369; // @[Main.scala 414:40 MemMap.scala 103:14]
  assign spriteRam_io_portA_wr = io_gameIndex == 4'h4 ? cs_5 & writeStrobe : _GEN_1370; // @[Main.scala 414:40 MemMap.scala 104:14]
  assign spriteRam_io_portA_addr = _GEN_1445[14:0];
  assign spriteRam_io_portA_mask = io_gameIndex == 4'h4 ? _mainRam_io_mask_T : _GEN_1309; // @[Main.scala 414:40 MemMap.scala 106:16]
  assign spriteRam_io_portA_din = io_gameIndex == 4'h4 ? cpu_io_dout : _GEN_1310; // @[Main.scala 414:40 MemMap.scala 107:15]
  assign spriteRam_io_portB_rd = io_gpuMem_sprite_vram_rd; // @[Main.scala 137:22]
  assign spriteRam_io_portB_addr = io_gpuMem_sprite_vram_addr; // @[Main.scala 137:22]
  assign vram8x8_0_clock = clock;
  assign vram8x8_0_io_clockB = io_videoClock; // @[Main.scala 148:19]
  assign vram8x8_0_io_portA_rd = io_gameIndex == 4'h4 ? cs_9 & readStrobe : _GEN_1321; // @[Main.scala 414:40 MemMap.scala 103:14]
  assign vram8x8_0_io_portA_wr = io_gameIndex == 4'h4 ? cs_9 & writeStrobe : _GEN_1322; // @[Main.scala 414:40 MemMap.scala 104:14]
  assign vram8x8_0_io_portA_addr = _GEN_1445[12:0];
  assign vram8x8_0_io_portA_mask = io_gameIndex == 4'h4 ? _mainRam_io_mask_T : _GEN_1309; // @[Main.scala 414:40 MemMap.scala 106:16]
  assign vram8x8_0_io_portA_din = io_gameIndex == 4'h4 ? cpu_io_dout : _GEN_1310; // @[Main.scala 414:40 MemMap.scala 107:15]
  assign vram8x8_0_io_portB_addr = io_gpuMem_layer_0_vram8x8_addr; // @[Main.scala 150:18]
  assign vram8x8_1_clock = clock;
  assign vram8x8_1_io_clockB = io_videoClock; // @[Main.scala 148:19]
  assign vram8x8_1_io_portA_rd = io_gameIndex == 4'h7 ? cs_194 & readStrobe : _GEN_1137; // @[Main.scala 393:42 MemMap.scala 103:14]
  assign vram8x8_1_io_portA_wr = io_gameIndex == 4'h7 ? cs_194 & writeStrobe : _GEN_1138; // @[Main.scala 393:42 MemMap.scala 104:14]
  assign vram8x8_1_io_portA_addr = _GEN_1308[12:0];
  assign vram8x8_1_io_portA_mask = io_gameIndex == 4'h7 ? _mainRam_io_mask_T : _GEN_1109; // @[Main.scala 393:42 MemMap.scala 106:16]
  assign vram8x8_1_io_portA_din = io_gameIndex == 4'h7 ? cpu_io_dout : _GEN_1110; // @[Main.scala 393:42 MemMap.scala 107:15]
  assign vram8x8_1_io_portB_addr = io_gpuMem_layer_1_vram8x8_addr; // @[Main.scala 150:18]
  assign vram8x8_2_clock = clock;
  assign vram8x8_2_io_clockB = io_videoClock; // @[Main.scala 148:19]
  assign vram8x8_2_io_portA_rd = io_gameIndex == 4'h7 ? cs_199 & readStrobe : _GEN_1148; // @[Main.scala 393:42 MemMap.scala 103:14]
  assign vram8x8_2_io_portA_wr = io_gameIndex == 4'h7 ? cs_199 & writeStrobe : _GEN_1149; // @[Main.scala 393:42 MemMap.scala 104:14]
  assign vram8x8_2_io_portA_addr = _GEN_1343[12:0];
  assign vram8x8_2_io_portA_mask = io_gameIndex == 4'h7 ? _mainRam_io_mask_T : _GEN_1151; // @[Main.scala 393:42 MemMap.scala 106:16]
  assign vram8x8_2_io_portA_din = io_gameIndex == 4'h7 ? cpu_io_dout : _GEN_1152; // @[Main.scala 393:42 MemMap.scala 107:15]
  assign vram8x8_2_io_portB_addr = io_gpuMem_layer_2_vram8x8_addr; // @[Main.scala 150:18]
  assign vram16x16_0_clock = clock;
  assign vram16x16_0_io_clockB = io_videoClock; // @[Main.scala 163:19]
  assign vram16x16_0_io_portA_rd = io_gameIndex == 4'h4 ? cs_6 & readStrobe : _GEN_1315; // @[Main.scala 414:40 MemMap.scala 103:14]
  assign vram16x16_0_io_portA_wr = io_gameIndex == 4'h4 ? cs_6 & writeStrobe : _GEN_1316; // @[Main.scala 414:40 MemMap.scala 104:14]
  assign vram16x16_0_io_portA_addr = _GEN_1445[10:0];
  assign vram16x16_0_io_portA_mask = io_gameIndex == 4'h4 ? _mainRam_io_mask_T : _GEN_1309; // @[Main.scala 414:40 MemMap.scala 106:16]
  assign vram16x16_0_io_portA_din = io_gameIndex == 4'h4 ? cpu_io_dout : _GEN_1310; // @[Main.scala 414:40 MemMap.scala 107:15]
  assign vram16x16_0_io_portB_addr = io_gpuMem_layer_0_vram16x16_addr; // @[Main.scala 165:18]
  assign vram16x16_1_clock = clock;
  assign vram16x16_1_io_clockB = io_videoClock; // @[Main.scala 163:19]
  assign vram16x16_1_io_portA_rd = io_gameIndex == 4'h7 ? cs_191 & readStrobe : _GEN_1131; // @[Main.scala 393:42 MemMap.scala 103:14]
  assign vram16x16_1_io_portA_wr = io_gameIndex == 4'h7 ? cs_191 & writeStrobe : _GEN_1132; // @[Main.scala 393:42 MemMap.scala 104:14]
  assign vram16x16_1_io_portA_addr = _GEN_1308[10:0];
  assign vram16x16_1_io_portA_mask = io_gameIndex == 4'h7 ? _mainRam_io_mask_T : _GEN_1109; // @[Main.scala 393:42 MemMap.scala 106:16]
  assign vram16x16_1_io_portA_din = io_gameIndex == 4'h7 ? cpu_io_dout : _GEN_1110; // @[Main.scala 393:42 MemMap.scala 107:15]
  assign vram16x16_1_io_portB_addr = io_gpuMem_layer_1_vram16x16_addr; // @[Main.scala 165:18]
  assign vram16x16_2_clock = clock;
  assign vram16x16_2_io_clockB = io_videoClock; // @[Main.scala 163:19]
  assign vram16x16_2_io_portA_rd = io_gameIndex == 4'h7 ? cs_196 & readStrobe : _GEN_1140; // @[Main.scala 393:42 MemMap.scala 103:14]
  assign vram16x16_2_io_portA_wr = io_gameIndex == 4'h7 ? cs_196 & writeStrobe : _GEN_1141; // @[Main.scala 393:42 MemMap.scala 104:14]
  assign vram16x16_2_io_portA_addr = _GEN_1335[10:0];
  assign vram16x16_2_io_portA_mask = io_gameIndex == 4'h7 ? _mainRam_io_mask_T : _GEN_1143; // @[Main.scala 393:42 MemMap.scala 106:16]
  assign vram16x16_2_io_portA_din = io_gameIndex == 4'h7 ? cpu_io_dout : _GEN_1144; // @[Main.scala 393:42 MemMap.scala 107:15]
  assign vram16x16_2_io_portB_addr = io_gpuMem_layer_2_vram16x16_addr; // @[Main.scala 165:18]
  assign lineRam_0_clock = clock;
  assign lineRam_0_io_clockB = io_videoClock; // @[Main.scala 178:19]
  assign lineRam_0_io_portA_rd = io_gameIndex == 4'h4 ? cs_7 & readStrobe : _GEN_1318; // @[Main.scala 414:40 MemMap.scala 103:14]
  assign lineRam_0_io_portA_wr = io_gameIndex == 4'h4 ? cs_7 & writeStrobe : _GEN_1319; // @[Main.scala 414:40 MemMap.scala 104:14]
  assign lineRam_0_io_portA_addr = _GEN_1445[9:0];
  assign lineRam_0_io_portA_mask = io_gameIndex == 4'h4 ? _mainRam_io_mask_T : _GEN_1309; // @[Main.scala 414:40 MemMap.scala 106:16]
  assign lineRam_0_io_portA_din = io_gameIndex == 4'h4 ? cpu_io_dout : _GEN_1310; // @[Main.scala 414:40 MemMap.scala 107:15]
  assign lineRam_0_io_portB_addr = io_gpuMem_layer_0_lineRam_addr; // @[Main.scala 180:18]
  assign lineRam_1_clock = clock;
  assign lineRam_1_io_clockB = io_videoClock; // @[Main.scala 178:19]
  assign lineRam_1_io_portA_rd = io_gameIndex == 4'h7 ? cs_192 & readStrobe : _GEN_1134; // @[Main.scala 393:42 MemMap.scala 103:14]
  assign lineRam_1_io_portA_wr = io_gameIndex == 4'h7 ? cs_192 & writeStrobe : _GEN_1135; // @[Main.scala 393:42 MemMap.scala 104:14]
  assign lineRam_1_io_portA_addr = _GEN_1308[9:0];
  assign lineRam_1_io_portA_mask = io_gameIndex == 4'h7 ? _mainRam_io_mask_T : _GEN_1109; // @[Main.scala 393:42 MemMap.scala 106:16]
  assign lineRam_1_io_portA_din = io_gameIndex == 4'h7 ? cpu_io_dout : _GEN_1110; // @[Main.scala 393:42 MemMap.scala 107:15]
  assign lineRam_1_io_portB_addr = io_gpuMem_layer_1_lineRam_addr; // @[Main.scala 180:18]
  assign lineRam_2_clock = clock;
  assign lineRam_2_io_clockB = io_videoClock; // @[Main.scala 178:19]
  assign lineRam_2_io_portA_rd = io_gameIndex == 4'h7 ? cs_197 & readStrobe : _GEN_1145; // @[Main.scala 393:42 MemMap.scala 103:14]
  assign lineRam_2_io_portA_wr = io_gameIndex == 4'h7 ? cs_197 & writeStrobe : _GEN_1146; // @[Main.scala 393:42 MemMap.scala 104:14]
  assign lineRam_2_io_portA_addr = _GEN_1335[9:0];
  assign lineRam_2_io_portA_mask = io_gameIndex == 4'h7 ? _mainRam_io_mask_T : _GEN_1143; // @[Main.scala 393:42 MemMap.scala 106:16]
  assign lineRam_2_io_portA_din = io_gameIndex == 4'h7 ? cpu_io_dout : _GEN_1144; // @[Main.scala 393:42 MemMap.scala 107:15]
  assign lineRam_2_io_portB_addr = io_gpuMem_layer_2_lineRam_addr; // @[Main.scala 180:18]
  assign paletteRam_clock = clock;
  assign paletteRam_io_clockB = io_videoClock; // @[Main.scala 192:24]
  assign paletteRam_io_portA_rd = io_gameIndex == 4'h4 ? cs_228 & readStrobe : _GEN_1311; // @[Main.scala 414:40 MemMap.scala 103:14]
  assign paletteRam_io_portA_wr = io_gameIndex == 4'h4 ? cs_228 & writeStrobe : _GEN_1312; // @[Main.scala 414:40 MemMap.scala 104:14]
  assign paletteRam_io_portA_addr = _GEN_1478[14:0];
  assign paletteRam_io_portA_mask = io_gameIndex == 4'h4 ? _mainRam_io_mask_T : _GEN_1309; // @[Main.scala 414:40 MemMap.scala 106:16]
  assign paletteRam_io_portA_din = io_gameIndex == 4'h4 ? cpu_io_dout : _GEN_1310; // @[Main.scala 414:40 MemMap.scala 107:15]
  assign paletteRam_io_portB_addr = io_gpuMem_paletteRam_addr; // @[Main.scala 194:23]
  assign layerRegs_0_clock = clock;
  assign layerRegs_0_io_mem_wr = io_gameIndex == 4'h4 ? cs_42 & writeStrobe : _GEN_1356; // @[Main.scala 414:40 MemMap.scala 104:14]
  assign layerRegs_0_io_mem_addr = _GEN_1445[1:0];
  assign layerRegs_0_io_mem_mask = io_gameIndex == 4'h4 ? _mainRam_io_mask_T : _GEN_1309; // @[Main.scala 414:40 MemMap.scala 106:16]
  assign layerRegs_0_io_mem_din = io_gameIndex == 4'h4 ? cpu_io_dout : _GEN_1310; // @[Main.scala 414:40 MemMap.scala 107:15]
  assign layerRegs_1_clock = clock;
  assign layerRegs_1_io_mem_wr = io_gameIndex == 4'h7 ? cs_207 & writeStrobe : _GEN_1162; // @[Main.scala 393:42 MemMap.scala 104:14]
  assign layerRegs_1_io_mem_addr = _GEN_1308[1:0];
  assign layerRegs_1_io_mem_mask = io_gameIndex == 4'h7 ? _mainRam_io_mask_T : _GEN_1109; // @[Main.scala 393:42 MemMap.scala 106:16]
  assign layerRegs_1_io_mem_din = io_gameIndex == 4'h7 ? cpu_io_dout : _GEN_1110; // @[Main.scala 393:42 MemMap.scala 107:15]
  assign layerRegs_2_clock = clock;
  assign layerRegs_2_io_mem_wr = io_gameIndex == 4'h7 ? cs_208 & writeStrobe : _GEN_1165; // @[Main.scala 393:42 MemMap.scala 104:14]
  assign layerRegs_2_io_mem_addr = _GEN_1363[1:0];
  assign layerRegs_2_io_mem_mask = io_gameIndex == 4'h7 ? _mainRam_io_mask_T : _GEN_1151; // @[Main.scala 393:42 MemMap.scala 106:16]
  assign layerRegs_2_io_mem_din = io_gameIndex == 4'h7 ? cpu_io_dout : _GEN_1152; // @[Main.scala 393:42 MemMap.scala 107:15]
  assign spriteRegs_clock = clock;
  assign spriteRegs_io_mem_wr = io_gameIndex == 4'h4 ? mem_7_wr : _GEN_1349; // @[Main.scala 414:40 MemIO.scala 305:8]
  assign spriteRegs_io_mem_addr = io_gameIndex == 4'h4 ? mem_addr : _GEN_1350; // @[Main.scala 414:40 MemIO.scala 306:10]
  assign spriteRegs_io_mem_mask = io_gameIndex == 4'h4 ? _mainRam_io_mask_T : _GEN_1309; // @[Main.scala 414:40 MemIO.scala 307:10]
  assign spriteRegs_io_mem_din = io_gameIndex == 4'h4 ? _GEN_193 : _GEN_1352; // @[Main.scala 414:40 MemIO.scala 308:9]
  always @(posedge clock) begin
    vBlank_r <= io_video_vBlank; // @[Reg.scala 19:16 20:{18,22}]
    vBlank <= vBlank_r; // @[Reg.scala 19:16 20:{18,22}]
    vBlankRising_REG <= vBlank; // @[Util.scala 158:44]
    pauseReg_REG <= io_player_0_pause | io_player_1_pause; // @[Main.scala 83:61]
    if (reset) begin // @[Util.scala 242:26]
      pauseReg <= 1'h0; // @[Util.scala 242:26]
    end else if (_pauseReg_T_2) begin // @[Util.scala 243:18]
      pauseReg <= ~pauseReg; // @[Util.scala 243:28]
    end
    if (reset) begin // @[Main.scala 86:25]
      videoIrq <= 1'h0; // @[Main.scala 86:25]
    end else if (io_gameIndex == 4'h4) begin // @[Main.scala 414:40]
      if (cs_223 & readStrobe) begin // @[MemMap.scala 180:30]
        if (offset_10 == 24'h4) begin // @[Main.scala 222:26]
          videoIrq <= 1'h0; // @[Main.scala 222:37]
        end else begin
          videoIrq <= _GEN_1346;
        end
      end else begin
        videoIrq <= _GEN_1346;
      end
    end else begin
      videoIrq <= _GEN_1346;
    end
    if (reset) begin // @[Main.scala 87:27]
      agalletIrq <= 1'h0; // @[Main.scala 87:27]
    end else begin
      agalletIrq <= _GEN_62;
    end
    if (reset) begin // @[MemMap.scala 48:23]
      dinReg <= 16'h0; // @[MemMap.scala 48:23]
    end else if (io_gameIndex == 4'h4) begin // @[Main.scala 414:40]
      if (cs_230 & readStrobe) begin // @[MemMap.scala 180:30]
        if (4'h5 == io_gameIndex) begin // @[Mux.scala 81:58]
          dinReg <= _right_T_9;
        end else begin
          dinReg <= _right_T_11;
        end
      end else if (cs_229 & readStrobe) begin // @[MemMap.scala 180:30]
        dinReg <= input0; // @[MemMap.scala 181:16]
      end else begin
        dinReg <= _GEN_1427;
      end
    end else if (io_gameIndex == 4'h7) begin // @[Main.scala 393:42]
      if (cs_213) begin // @[MemMap.scala 108:16]
        dinReg <= spriteRam_io_portA_dout; // @[MemMap.scala 109:16]
      end else begin
        dinReg <= _GEN_1295;
      end
    end else if (_cs_T) begin // @[Main.scala 368:41]
      dinReg <= _GEN_1098;
    end else begin
      dinReg <= _GEN_897;
    end
    if (reset) begin // @[MemMap.scala 49:25]
      dtackReg <= 1'h0; // @[MemMap.scala 49:25]
    end else if (io_gameIndex == 4'h4) begin // @[Main.scala 414:40]
      dtackReg <= _GEN_1436;
    end else if (io_gameIndex == 4'h7) begin // @[Main.scala 393:42]
      dtackReg <= _GEN_1299;
    end else if (_cs_T) begin // @[Main.scala 368:41]
      dtackReg <= _GEN_1099;
    end else begin
      dtackReg <= _GEN_892;
    end
    readStrobe_REG <= cpu_io_as; // @[Util.scala 158:44]
    upperWriteStrobe_REG <= cpu_io_uds; // @[Util.scala 158:44]
    lowerWriteStrobe_REG <= cpu_io_lds; // @[Util.scala 158:44]
    if (reset) begin // @[Reg.scala 35:20]
      eeprom_io_serial_cs_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (eepromMem_wr) begin // @[Reg.scala 36:18]
      if (io_gameIndex == 4'h5) begin // @[Main.scala 111:15]
        eeprom_io_serial_cs_r <= eepromMem_din[5];
      end else begin
        eeprom_io_serial_cs_r <= eepromMem_din[9];
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      eeprom_io_serial_sck_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (eepromMem_wr) begin // @[Reg.scala 36:18]
      if (_cs_T) begin // @[Main.scala 112:16]
        eeprom_io_serial_sck_r <= eepromMem_din[6];
      end else begin
        eeprom_io_serial_sck_r <= eepromMem_din[10];
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      eeprom_io_serial_sdi_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (eepromMem_wr) begin // @[Reg.scala 36:18]
      if (_cs_T) begin // @[Main.scala 113:16]
        eeprom_io_serial_sdi_r <= eepromMem_din[7];
      end else begin
        eeprom_io_serial_sdi_r <= eepromMem_din[11];
      end
    end
    REG <= vBlank; // @[Util.scala 165:45]
    if (reset) begin // @[Counter.scala 40:34]
      coin1_pulseCounterWrap_value <= 22'h0; // @[Counter.scala 40:34]
    end else if (coin1_s_enableReg) begin // @[Counter.scala 86:48]
      if (coin1_pulseCounterWrap_wrap_wrap) begin // @[Counter.scala 48:20]
        coin1_pulseCounterWrap_value <= 22'h0; // @[Counter.scala 48:28]
      end else begin
        coin1_pulseCounterWrap_value <= _coin1_pulseCounterWrap_wrap_value_T_1; // @[Counter.scala 46:13]
      end
    end
    if (reset) begin // @[Util.scala 218:28]
      coin1_s_enableReg <= 1'h0; // @[Util.scala 218:28]
    end else if (coin1_pulseCounterWrap) begin // @[Util.scala 219:17]
      coin1_s_enableReg <= 1'h0; // @[Util.scala 219:29]
    end else begin
      coin1_s_enableReg <= _GEN_68;
    end
    coin1_s_REG <= io_player_0_coin; // @[Util.scala 158:44]
    if (reset) begin // @[Counter.scala 40:34]
      coin2_pulseCounterWrap_value <= 22'h0; // @[Counter.scala 40:34]
    end else if (coin2_s_enableReg) begin // @[Counter.scala 86:48]
      if (coin2_pulseCounterWrap_wrap_wrap) begin // @[Counter.scala 48:20]
        coin2_pulseCounterWrap_value <= 22'h0; // @[Counter.scala 48:28]
      end else begin
        coin2_pulseCounterWrap_value <= _coin2_pulseCounterWrap_wrap_value_T_1; // @[Counter.scala 46:13]
      end
    end
    if (reset) begin // @[Util.scala 218:28]
      coin2_s_enableReg <= 1'h0; // @[Util.scala 218:28]
    end else if (coin2_pulseCounterWrap) begin // @[Util.scala 219:17]
      coin2_s_enableReg <= 1'h0; // @[Util.scala 219:29]
    end else begin
      coin2_s_enableReg <= _GEN_75;
    end
    coin2_s_REG <= io_player_1_coin; // @[Util.scala 158:44]
    if (reset) begin // @[Counter.scala 40:34]
      service_pulseCounterWrap_value <= 27'h0; // @[Counter.scala 40:34]
    end else if (service_s_enableReg) begin // @[Counter.scala 86:48]
      if (service_pulseCounterWrap_wrap_wrap) begin // @[Counter.scala 48:20]
        service_pulseCounterWrap_value <= 27'h0; // @[Counter.scala 48:28]
      end else begin
        service_pulseCounterWrap_value <= _service_pulseCounterWrap_wrap_value_T_1; // @[Counter.scala 46:13]
      end
    end
    if (reset) begin // @[Util.scala 218:28]
      service_s_enableReg <= 1'h0; // @[Util.scala 218:28]
    end else if (service_pulseCounterWrap) begin // @[Util.scala 219:17]
      service_s_enableReg <= 1'h0; // @[Util.scala 219:29]
    end else begin
      service_s_enableReg <= _GEN_82;
    end
    service_s_REG <= io_options_service; // @[Util.scala 158:44]
    if (cs_8) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_10) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_1 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_13) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_2 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_15) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_3 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_31) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_4 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_33) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_5 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_36) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_6 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_38) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_7 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_8) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_8 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_10) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_9 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_13) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_10 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_15) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_11 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_8) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_12 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_10) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_13 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_13) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_14 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_15) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_15 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_98) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_16 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_100) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_17 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_8) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_18 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_10) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_19 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_13) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_20 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_15) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_21 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_98) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_22 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_100) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_23 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_8) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_24 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_10) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_25 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_13) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_26 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_15) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_27 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_98) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_28 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_100) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_29 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_188) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_30 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_190) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_31 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_193) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_32 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_195) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_33 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_198) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_34 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_200) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_35 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_8) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_36 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
    if (cs_10) begin // @[MemMap.scala 164:16]
      if (!(readStrobe)) begin // @[MemMap.scala 165:26]
        if (writeStrobe) begin // @[MemMap.scala 167:33]
          tmp_37 <= cpu_io_dout; // @[MemMap.scala 207:45]
        end
      end
    end
  end
  always @(posedge io_videoClock) begin
    io_gpuMem_layer_0_regs_r_tileSize <= layerRegs_0_io_regs_1[13]; // @[LayerRegs.scala 83:29]
    io_gpuMem_layer_0_regs_r_enable <= ~layerRegs_0_io_regs_2[4]; // @[LayerRegs.scala 84:20]
    io_gpuMem_layer_0_regs_r_flipX <= ~layerRegs_0_io_regs_0[15]; // @[LayerRegs.scala 85:19]
    io_gpuMem_layer_0_regs_r_flipY <= ~layerRegs_0_io_regs_1[15]; // @[LayerRegs.scala 86:19]
    io_gpuMem_layer_0_regs_r_rowScrollEnable <= layerRegs_0_io_regs_0[14]; // @[LayerRegs.scala 87:36]
    io_gpuMem_layer_0_regs_r_rowSelectEnable <= layerRegs_0_io_regs_1[14]; // @[LayerRegs.scala 88:36]
    io_gpuMem_layer_0_regs_r_scroll_x <= layerRegs_0_io_regs_0[8:0]; // @[LayerRegs.scala 89:33]
    io_gpuMem_layer_0_regs_r_scroll_y <= layerRegs_0_io_regs_1[8:0]; // @[LayerRegs.scala 89:48]
    io_gpuMem_layer_0_regs_r_1_tileSize <= io_gpuMem_layer_0_regs_r_tileSize; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_0_regs_r_1_enable <= io_gpuMem_layer_0_regs_r_enable; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_0_regs_r_1_flipX <= io_gpuMem_layer_0_regs_r_flipX; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_0_regs_r_1_flipY <= io_gpuMem_layer_0_regs_r_flipY; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_0_regs_r_1_rowScrollEnable <= io_gpuMem_layer_0_regs_r_rowScrollEnable; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_0_regs_r_1_rowSelectEnable <= io_gpuMem_layer_0_regs_r_rowSelectEnable; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_0_regs_r_1_scroll_x <= io_gpuMem_layer_0_regs_r_scroll_x; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_0_regs_r_1_scroll_y <= io_gpuMem_layer_0_regs_r_scroll_y; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_1_regs_r_tileSize <= layerRegs_1_io_regs_1[13]; // @[LayerRegs.scala 83:29]
    io_gpuMem_layer_1_regs_r_enable <= ~layerRegs_1_io_regs_2[4]; // @[LayerRegs.scala 84:20]
    io_gpuMem_layer_1_regs_r_flipX <= ~layerRegs_1_io_regs_0[15]; // @[LayerRegs.scala 85:19]
    io_gpuMem_layer_1_regs_r_flipY <= ~layerRegs_1_io_regs_1[15]; // @[LayerRegs.scala 86:19]
    io_gpuMem_layer_1_regs_r_rowScrollEnable <= layerRegs_1_io_regs_0[14]; // @[LayerRegs.scala 87:36]
    io_gpuMem_layer_1_regs_r_rowSelectEnable <= layerRegs_1_io_regs_1[14]; // @[LayerRegs.scala 88:36]
    io_gpuMem_layer_1_regs_r_scroll_x <= layerRegs_1_io_regs_0[8:0]; // @[LayerRegs.scala 89:33]
    io_gpuMem_layer_1_regs_r_scroll_y <= layerRegs_1_io_regs_1[8:0]; // @[LayerRegs.scala 89:48]
    io_gpuMem_layer_1_regs_r_1_tileSize <= io_gpuMem_layer_1_regs_r_tileSize; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_1_regs_r_1_enable <= io_gpuMem_layer_1_regs_r_enable; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_1_regs_r_1_flipX <= io_gpuMem_layer_1_regs_r_flipX; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_1_regs_r_1_flipY <= io_gpuMem_layer_1_regs_r_flipY; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_1_regs_r_1_rowScrollEnable <= io_gpuMem_layer_1_regs_r_rowScrollEnable; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_1_regs_r_1_rowSelectEnable <= io_gpuMem_layer_1_regs_r_rowSelectEnable; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_1_regs_r_1_scroll_x <= io_gpuMem_layer_1_regs_r_scroll_x; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_1_regs_r_1_scroll_y <= io_gpuMem_layer_1_regs_r_scroll_y; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_2_regs_r_tileSize <= layerRegs_2_io_regs_1[13]; // @[LayerRegs.scala 83:29]
    io_gpuMem_layer_2_regs_r_enable <= ~layerRegs_2_io_regs_2[4]; // @[LayerRegs.scala 84:20]
    io_gpuMem_layer_2_regs_r_flipX <= ~layerRegs_2_io_regs_0[15]; // @[LayerRegs.scala 85:19]
    io_gpuMem_layer_2_regs_r_flipY <= ~layerRegs_2_io_regs_1[15]; // @[LayerRegs.scala 86:19]
    io_gpuMem_layer_2_regs_r_rowScrollEnable <= layerRegs_2_io_regs_0[14]; // @[LayerRegs.scala 87:36]
    io_gpuMem_layer_2_regs_r_rowSelectEnable <= layerRegs_2_io_regs_1[14]; // @[LayerRegs.scala 88:36]
    io_gpuMem_layer_2_regs_r_scroll_x <= layerRegs_2_io_regs_0[8:0]; // @[LayerRegs.scala 89:33]
    io_gpuMem_layer_2_regs_r_scroll_y <= layerRegs_2_io_regs_1[8:0]; // @[LayerRegs.scala 89:48]
    io_gpuMem_layer_2_regs_r_1_tileSize <= io_gpuMem_layer_2_regs_r_tileSize; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_2_regs_r_1_enable <= io_gpuMem_layer_2_regs_r_enable; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_2_regs_r_1_flipX <= io_gpuMem_layer_2_regs_r_flipX; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_2_regs_r_1_flipY <= io_gpuMem_layer_2_regs_r_flipY; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_2_regs_r_1_rowScrollEnable <= io_gpuMem_layer_2_regs_r_rowScrollEnable; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_2_regs_r_1_rowSelectEnable <= io_gpuMem_layer_2_regs_r_rowSelectEnable; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_2_regs_r_1_scroll_x <= io_gpuMem_layer_2_regs_r_scroll_x; // @[Reg.scala 19:16 20:{18,22}]
    io_gpuMem_layer_2_regs_r_1_scroll_y <= io_gpuMem_layer_2_regs_r_scroll_y; // @[Reg.scala 19:16 20:{18,22}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  vBlank_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  vBlank = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  vBlankRising_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pauseReg_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pauseReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  videoIrq = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  agalletIrq = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dinReg = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  dtackReg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  readStrobe_REG = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  upperWriteStrobe_REG = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  lowerWriteStrobe_REG = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  eeprom_io_serial_cs_r = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  eeprom_io_serial_sck_r = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  eeprom_io_serial_sdi_r = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_tileSize = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_enable = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_flipX = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_flipY = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_rowScrollEnable = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_rowSelectEnable = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_scroll_x = _RAND_21[8:0];
  _RAND_22 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_scroll_y = _RAND_22[8:0];
  _RAND_23 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_1_tileSize = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_1_enable = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_1_flipX = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_1_flipY = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_1_rowScrollEnable = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_1_rowSelectEnable = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_1_scroll_x = _RAND_29[8:0];
  _RAND_30 = {1{`RANDOM}};
  io_gpuMem_layer_0_regs_r_1_scroll_y = _RAND_30[8:0];
  _RAND_31 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_tileSize = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_enable = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_flipX = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_flipY = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_rowScrollEnable = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_rowSelectEnable = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_scroll_x = _RAND_37[8:0];
  _RAND_38 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_scroll_y = _RAND_38[8:0];
  _RAND_39 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_1_tileSize = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_1_enable = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_1_flipX = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_1_flipY = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_1_rowScrollEnable = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_1_rowSelectEnable = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_1_scroll_x = _RAND_45[8:0];
  _RAND_46 = {1{`RANDOM}};
  io_gpuMem_layer_1_regs_r_1_scroll_y = _RAND_46[8:0];
  _RAND_47 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_tileSize = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_enable = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_flipX = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_flipY = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_rowScrollEnable = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_rowSelectEnable = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_scroll_x = _RAND_53[8:0];
  _RAND_54 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_scroll_y = _RAND_54[8:0];
  _RAND_55 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_1_tileSize = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_1_enable = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_1_flipX = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_1_flipY = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_1_rowScrollEnable = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_1_rowSelectEnable = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_1_scroll_x = _RAND_61[8:0];
  _RAND_62 = {1{`RANDOM}};
  io_gpuMem_layer_2_regs_r_1_scroll_y = _RAND_62[8:0];
  _RAND_63 = {1{`RANDOM}};
  REG = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  coin1_pulseCounterWrap_value = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  coin1_s_enableReg = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  coin1_s_REG = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  coin2_pulseCounterWrap_value = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  coin2_s_enableReg = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  coin2_s_REG = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  service_pulseCounterWrap_value = _RAND_70[26:0];
  _RAND_71 = {1{`RANDOM}};
  service_s_enableReg = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  service_s_REG = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  tmp = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  tmp_1 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  tmp_2 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  tmp_3 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  tmp_4 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  tmp_5 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  tmp_6 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  tmp_7 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  tmp_8 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  tmp_9 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  tmp_10 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  tmp_11 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  tmp_12 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  tmp_13 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  tmp_14 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  tmp_15 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  tmp_16 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  tmp_17 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  tmp_18 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  tmp_19 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  tmp_20 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  tmp_21 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  tmp_22 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  tmp_23 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  tmp_24 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  tmp_25 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  tmp_26 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  tmp_27 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  tmp_28 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  tmp_29 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  tmp_30 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  tmp_31 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  tmp_32 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  tmp_33 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  tmp_34 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  tmp_35 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  tmp_36 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  tmp_37 = _RAND_110[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReadDataFreezer(
  input         clock,
  input         reset,
  input         io_targetClock,
  input         io_in_rd,
  input  [19:0] io_in_addr,
  output [15:0] io_in_dout,
  output        io_in_valid,
  output        io_out_rd,
  output [19:0] io_out_addr,
  input  [15:0] io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg  clear_s; // @[Util.scala 242:26]
  wire  _clear_s_dataReg_T = ~clear_s; // @[Util.scala 243:31]
  reg  clear_REG; // @[Util.scala 151:40]
  wire  clear = clear_s ^ clear_REG; // @[Util.scala 151:31]
  wire  _wait_n_T = ~clear; // @[Util.scala 190:24]
  reg  valid_enableReg; // @[Util.scala 188:28]
  wire  _GEN_3 = clear ? 1'h0 : valid_enableReg; // @[Util.scala 188:28 189:{53,65}]
  wire  _GEN_4 = io_out_valid | _GEN_3; // @[Util.scala 189:{13,25}]
  reg [15:0] data_dataReg; // @[Reg.scala 19:16]
  reg  data_enableReg; // @[Util.scala 204:28]
  wire  _GEN_6 = io_out_valid | data_enableReg; // @[Util.scala 204:28 205:{54,66}]
  reg  pendingRead; // @[Crossing.scala 116:28]
  wire  effectiveRead = io_in_rd & io_out_wait_n; // @[Crossing.scala 117:32]
  reg  clearRead_REG; // @[Crossing.scala 118:35]
  wire  clearRead = clear & clearRead_REG; // @[Crossing.scala 118:25]
  wire  _GEN_8 = clearRead ? 1'h0 : pendingRead; // @[Crossing.scala 116:28 119:{69,83}]
  wire  _GEN_9 = effectiveRead | _GEN_8; // @[Crossing.scala 119:{23,37}]
  assign io_in_dout = data_enableReg & _wait_n_T ? data_dataReg : io_out_dout; // @[Util.scala 206:8]
  assign io_in_valid = io_out_valid | valid_enableReg & ~clear; // @[Util.scala 190:7]
  assign io_out_rd = io_in_rd & (~pendingRead | clearRead); // @[Crossing.scala 128:25]
  assign io_out_addr = io_in_addr; // @[Crossing.scala 122:9]
  always @(posedge io_targetClock) begin
    if (reset) begin // @[Util.scala 242:26]
      clear_s <= 1'h0; // @[Util.scala 242:26]
    end else begin
      clear_s <= _clear_s_dataReg_T;
    end
  end
  always @(posedge clock) begin
    clear_REG <= clear_s; // @[Util.scala 151:40]
    if (reset) begin // @[Util.scala 188:28]
      valid_enableReg <= 1'h0; // @[Util.scala 188:28]
    end else begin
      valid_enableReg <= _GEN_4;
    end
    if (io_out_valid) begin // @[Reg.scala 20:18]
      data_dataReg <= io_out_dout; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[Util.scala 204:28]
      data_enableReg <= 1'h0; // @[Util.scala 204:28]
    end else if (clear) begin // @[Util.scala 205:17]
      data_enableReg <= 1'h0; // @[Util.scala 205:29]
    end else begin
      data_enableReg <= _GEN_6;
    end
    if (reset) begin // @[Crossing.scala 116:28]
      pendingRead <= 1'h0; // @[Crossing.scala 116:28]
    end else begin
      pendingRead <= _GEN_9;
    end
    clearRead_REG <= io_out_valid | valid_enableReg & ~clear; // @[Util.scala 190:7]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  clear_s = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  clear_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  valid_enableReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  data_dataReg = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  data_enableReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  pendingRead = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  clearRead_REG = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DataFreezer(
  input         clock,
  input         reset,
  input         io_targetClock,
  input         io_in_rd,
  input         io_in_wr,
  input  [6:0]  io_in_addr,
  input  [15:0] io_in_din,
  output [15:0] io_in_dout,
  output        io_in_wait_n,
  output        io_in_valid,
  output        io_out_rd,
  output        io_out_wr,
  output [6:0]  io_out_addr,
  output [15:0] io_out_din,
  input  [15:0] io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  clear_s; // @[Util.scala 242:26]
  wire  _clear_s_dataReg_T = ~clear_s; // @[Util.scala 243:31]
  reg  clear_REG; // @[Util.scala 151:40]
  wire  clear = clear_s ^ clear_REG; // @[Util.scala 151:31]
  reg  wait_n_enableReg; // @[Util.scala 188:28]
  wire  _GEN_1 = clear ? 1'h0 : wait_n_enableReg; // @[Util.scala 188:28 189:{53,65}]
  wire  _GEN_2 = io_out_wait_n | _GEN_1; // @[Util.scala 189:{13,25}]
  wire  _wait_n_T = ~clear; // @[Util.scala 190:24]
  wire  wait_n = io_out_wait_n | wait_n_enableReg & ~clear; // @[Util.scala 190:7]
  reg  valid_enableReg; // @[Util.scala 188:28]
  wire  _GEN_3 = clear ? 1'h0 : valid_enableReg; // @[Util.scala 188:28 189:{53,65}]
  wire  _GEN_4 = io_out_valid | _GEN_3; // @[Util.scala 189:{13,25}]
  wire  valid = io_out_valid | valid_enableReg & ~clear; // @[Util.scala 190:7]
  reg [15:0] data_dataReg; // @[Reg.scala 19:16]
  reg  data_enableReg; // @[Util.scala 204:28]
  wire  _GEN_6 = io_out_valid | data_enableReg; // @[Util.scala 204:28 205:{54,66}]
  reg  pendingRead; // @[Crossing.scala 170:28]
  reg  pendingWrite; // @[Crossing.scala 171:29]
  wire  effectiveRead = io_in_rd & io_out_wait_n; // @[Crossing.scala 172:32]
  wire  effectiveWrite = io_in_wr & io_out_wait_n; // @[Crossing.scala 173:33]
  reg  clearRead_REG; // @[Crossing.scala 174:35]
  wire  clearRead = clear & clearRead_REG; // @[Crossing.scala 174:25]
  wire  _GEN_8 = clearRead ? 1'h0 : pendingRead; // @[Crossing.scala 170:28 176:{69,83}]
  wire  _GEN_9 = effectiveRead | _GEN_8; // @[Crossing.scala 176:{23,37}]
  wire  _GEN_10 = clear ? 1'h0 : pendingWrite; // @[Crossing.scala 171:29 177:{72,87}]
  wire  _GEN_11 = effectiveWrite | _GEN_10; // @[Crossing.scala 177:{24,39}]
  assign io_in_dout = data_enableReg & _wait_n_T ? data_dataReg : io_out_dout; // @[Util.scala 206:8]
  assign io_in_wait_n = io_out_wait_n | wait_n_enableReg & ~clear; // @[Util.scala 190:7]
  assign io_in_valid = io_out_valid | valid_enableReg & ~clear; // @[Util.scala 190:7]
  assign io_out_rd = io_in_rd & (~pendingRead | clearRead); // @[Crossing.scala 186:25]
  assign io_out_wr = io_in_wr & (~pendingWrite | clear); // @[Crossing.scala 187:25]
  assign io_out_addr = io_in_addr; // @[Crossing.scala 180:9]
  assign io_out_din = io_in_din; // @[Crossing.scala 180:9]
  always @(posedge io_targetClock) begin
    if (reset) begin // @[Util.scala 242:26]
      clear_s <= 1'h0; // @[Util.scala 242:26]
    end else begin
      clear_s <= _clear_s_dataReg_T;
    end
  end
  always @(posedge clock) begin
    clear_REG <= clear_s; // @[Util.scala 151:40]
    if (reset) begin // @[Util.scala 188:28]
      wait_n_enableReg <= 1'h0; // @[Util.scala 188:28]
    end else begin
      wait_n_enableReg <= _GEN_2;
    end
    if (reset) begin // @[Util.scala 188:28]
      valid_enableReg <= 1'h0; // @[Util.scala 188:28]
    end else begin
      valid_enableReg <= _GEN_4;
    end
    if (io_out_valid) begin // @[Reg.scala 20:18]
      data_dataReg <= io_out_dout; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[Util.scala 204:28]
      data_enableReg <= 1'h0; // @[Util.scala 204:28]
    end else if (clear) begin // @[Util.scala 205:17]
      data_enableReg <= 1'h0; // @[Util.scala 205:29]
    end else begin
      data_enableReg <= _GEN_6;
    end
    if (reset) begin // @[Crossing.scala 170:28]
      pendingRead <= 1'h0; // @[Crossing.scala 170:28]
    end else begin
      pendingRead <= _GEN_9;
    end
    if (reset) begin // @[Crossing.scala 171:29]
      pendingWrite <= 1'h0; // @[Crossing.scala 171:29]
    end else begin
      pendingWrite <= _GEN_11;
    end
    clearRead_REG <= io_out_valid | valid_enableReg & ~clear; // @[Util.scala 190:7]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"DataFreezer(read: %d, write: %d, wait: %d, valid: %d, clear: %d)\n",io_out_rd,io_out_wr,
            wait_n,valid,clear); // @[Crossing.scala 189:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  clear_s = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  clear_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wait_n_enableReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  valid_enableReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  data_dataReg = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  data_enableReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pendingRead = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pendingWrite = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  clearRead_REG = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CPU_1(
  input         clock,
  input         reset,
  output [15:0] io_addr,
  input  [7:0]  io_din,
  output [7:0]  io_dout,
  output        io_rd,
  output        io_wr,
  output        io_rfsh,
  output        io_mreq,
  output        io_iorq,
  input         io_int,
  input         io_nmi
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  cpu_RESET_n; // @[CPU.scala 101:19]
  wire  cpu_CLK; // @[CPU.scala 101:19]
  wire  cpu_CEN; // @[CPU.scala 101:19]
  wire  cpu_WAIT_n; // @[CPU.scala 101:19]
  wire  cpu_INT_n; // @[CPU.scala 101:19]
  wire  cpu_NMI_n; // @[CPU.scala 101:19]
  wire  cpu_BUSRQ_n; // @[CPU.scala 101:19]
  wire  cpu_M1_n; // @[CPU.scala 101:19]
  wire  cpu_MREQ_n; // @[CPU.scala 101:19]
  wire  cpu_IORQ_n; // @[CPU.scala 101:19]
  wire  cpu_RD_n; // @[CPU.scala 101:19]
  wire  cpu_WR_n; // @[CPU.scala 101:19]
  wire  cpu_RFSH_n; // @[CPU.scala 101:19]
  wire  cpu_HALT_n; // @[CPU.scala 101:19]
  wire  cpu_BUSAK_n; // @[CPU.scala 101:19]
  wire [15:0] cpu_A; // @[CPU.scala 101:19]
  wire [7:0] cpu_DI; // @[CPU.scala 101:19]
  wire [7:0] cpu_DO; // @[CPU.scala 101:19]
  wire [210:0] cpu_REG; // @[CPU.scala 101:19]
  reg [2:0] cen_value; // @[Counter.scala 40:34]
  wire [2:0] _cen_wrap_value_T_1 = cen_value + 3'h1; // @[Counter.scala 46:22]
  T80s cpu ( // @[CPU.scala 101:19]
    .RESET_n(cpu_RESET_n),
    .CLK(cpu_CLK),
    .CEN(cpu_CEN),
    .WAIT_n(cpu_WAIT_n),
    .INT_n(cpu_INT_n),
    .NMI_n(cpu_NMI_n),
    .BUSRQ_n(cpu_BUSRQ_n),
    .M1_n(cpu_M1_n),
    .MREQ_n(cpu_MREQ_n),
    .IORQ_n(cpu_IORQ_n),
    .RD_n(cpu_RD_n),
    .WR_n(cpu_WR_n),
    .RFSH_n(cpu_RFSH_n),
    .HALT_n(cpu_HALT_n),
    .BUSAK_n(cpu_BUSAK_n),
    .A(cpu_A),
    .DI(cpu_DI),
    .DO(cpu_DO),
    .REG(cpu_REG)
  );
  assign io_addr = cpu_A; // @[CPU.scala 117:11]
  assign io_dout = cpu_DO; // @[CPU.scala 118:11]
  assign io_rd = ~cpu_RD_n; // @[CPU.scala 112:12]
  assign io_wr = ~cpu_WR_n; // @[CPU.scala 113:12]
  assign io_rfsh = ~cpu_RFSH_n; // @[CPU.scala 114:14]
  assign io_mreq = ~cpu_MREQ_n; // @[CPU.scala 110:14]
  assign io_iorq = ~cpu_IORQ_n; // @[CPU.scala 111:14]
  assign cpu_RESET_n = ~reset; // @[CPU.scala 102:21]
  assign cpu_CLK = clock; // @[CPU.scala 103:14]
  assign cpu_CEN = cen_value == 3'h7; // @[Counter.scala 45:24]
  assign cpu_WAIT_n = 1'h1; // @[CPU.scala 105:20]
  assign cpu_INT_n = ~io_int; // @[CPU.scala 106:19]
  assign cpu_NMI_n = ~io_nmi; // @[CPU.scala 107:19]
  assign cpu_BUSRQ_n = 1'h1; // @[CPU.scala 108:18]
  assign cpu_DI = io_din; // @[CPU.scala 109:13]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 40:34]
      cen_value <= 3'h0; // @[Counter.scala 40:34]
    end else begin
      cen_value <= _cen_wrap_value_T_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cen_value = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SinglePortRam_1(
  input         clock,
  input         io_rd,
  input         io_wr,
  input  [12:0] io_addr,
  input  [7:0]  io_din,
  output [7:0]  io_dout
);
  wire  ram_clk; // @[SinglePortRam.scala 72:19]
  wire  ram_rd; // @[SinglePortRam.scala 72:19]
  wire  ram_wr; // @[SinglePortRam.scala 72:19]
  wire [12:0] ram_addr; // @[SinglePortRam.scala 72:19]
  wire  ram_mask; // @[SinglePortRam.scala 72:19]
  wire [7:0] ram_din; // @[SinglePortRam.scala 72:19]
  wire [7:0] ram_dout; // @[SinglePortRam.scala 72:19]
  single_port_ram #(.ADDR_WIDTH(13), .DATA_WIDTH(8), .DEPTH(0), .MASK_ENABLE("FALSE")) ram ( // @[SinglePortRam.scala 72:19]
    .clk(ram_clk),
    .rd(ram_rd),
    .wr(ram_wr),
    .addr(ram_addr),
    .mask(ram_mask),
    .din(ram_din),
    .dout(ram_dout)
  );
  assign io_dout = ram_dout; // @[SinglePortRam.scala 79:11]
  assign ram_clk = clock; // @[SinglePortRam.scala 73:14]
  assign ram_rd = io_rd; // @[SinglePortRam.scala 74:13]
  assign ram_wr = io_wr; // @[SinglePortRam.scala 75:13]
  assign ram_addr = io_addr; // @[SinglePortRam.scala 76:15]
  assign ram_mask = 1'h0; // @[SinglePortRam.scala 77:15]
  assign ram_din = io_din; // @[SinglePortRam.scala 78:14]
endmodule
module NMK112(
  input         clock,
  input         io_cpu_wr,
  input  [22:0] io_cpu_addr,
  input  [15:0] io_cpu_din,
  input  [24:0] io_addr_0_in,
  output [24:0] io_addr_0_out,
  input  [24:0] io_addr_1_in,
  output [24:0] io_addr_1_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] pageTableReg_0_0; // @[NMK112.scala 85:25]
  reg [4:0] pageTableReg_0_1; // @[NMK112.scala 85:25]
  reg [4:0] pageTableReg_0_2; // @[NMK112.scala 85:25]
  reg [4:0] pageTableReg_0_3; // @[NMK112.scala 85:25]
  reg [4:0] pageTableReg_1_0; // @[NMK112.scala 85:25]
  reg [4:0] pageTableReg_1_1; // @[NMK112.scala 85:25]
  reg [4:0] pageTableReg_1_2; // @[NMK112.scala 85:25]
  reg [4:0] pageTableReg_1_3; // @[NMK112.scala 85:25]
  wire  chip = io_cpu_addr[2]; // @[NMK112.scala 89:27]
  wire [1:0] bank = io_cpu_addr[1:0]; // @[NMK112.scala 90:27]
  wire [1:0] io_addr_0_out_bank = io_addr_0_in[17:16]; // @[NMK112.scala 127:48]
  wire [4:0] _GEN_17 = 2'h1 == io_addr_0_out_bank ? pageTableReg_0_1 : pageTableReg_0_0; // @[NMK112.scala 128:{21,21}]
  wire [4:0] _GEN_18 = 2'h2 == io_addr_0_out_bank ? pageTableReg_0_2 : _GEN_17; // @[NMK112.scala 128:{21,21}]
  wire [4:0] _GEN_19 = 2'h3 == io_addr_0_out_bank ? pageTableReg_0_3 : _GEN_18; // @[NMK112.scala 128:{21,21}]
  wire [20:0] _io_addr_0_out_T_2 = {_GEN_19,io_addr_0_in[15:0]}; // @[NMK112.scala 128:21]
  wire [1:0] io_addr_1_out_bank = io_addr_1_in > 25'h400 ? io_addr_1_in[17:16] : io_addr_1_in[9:8]; // @[NMK112.scala 127:19]
  wire [4:0] _GEN_21 = 2'h1 == io_addr_1_out_bank ? pageTableReg_1_1 : pageTableReg_1_0; // @[NMK112.scala 128:{21,21}]
  wire [4:0] _GEN_22 = 2'h2 == io_addr_1_out_bank ? pageTableReg_1_2 : _GEN_21; // @[NMK112.scala 128:{21,21}]
  wire [4:0] _GEN_23 = 2'h3 == io_addr_1_out_bank ? pageTableReg_1_3 : _GEN_22; // @[NMK112.scala 128:{21,21}]
  wire [20:0] _io_addr_1_out_T_2 = {_GEN_23,io_addr_1_in[15:0]}; // @[NMK112.scala 128:21]
  assign io_addr_0_out = {{4'd0}, _io_addr_0_out_T_2}; // @[NMK112.scala 96:20]
  assign io_addr_1_out = {{4'd0}, _io_addr_1_out_T_2}; // @[NMK112.scala 96:20]
  always @(posedge clock) begin
    if (io_cpu_wr) begin // @[NMK112.scala 88:19]
      if (~chip & 2'h0 == bank) begin // @[NMK112.scala 91:30]
        pageTableReg_0_0 <= io_cpu_din[4:0]; // @[NMK112.scala 91:30]
      end
    end
    if (io_cpu_wr) begin // @[NMK112.scala 88:19]
      if (~chip & 2'h1 == bank) begin // @[NMK112.scala 91:30]
        pageTableReg_0_1 <= io_cpu_din[4:0]; // @[NMK112.scala 91:30]
      end
    end
    if (io_cpu_wr) begin // @[NMK112.scala 88:19]
      if (~chip & 2'h2 == bank) begin // @[NMK112.scala 91:30]
        pageTableReg_0_2 <= io_cpu_din[4:0]; // @[NMK112.scala 91:30]
      end
    end
    if (io_cpu_wr) begin // @[NMK112.scala 88:19]
      if (~chip & 2'h3 == bank) begin // @[NMK112.scala 91:30]
        pageTableReg_0_3 <= io_cpu_din[4:0]; // @[NMK112.scala 91:30]
      end
    end
    if (io_cpu_wr) begin // @[NMK112.scala 88:19]
      if (chip & 2'h0 == bank) begin // @[NMK112.scala 91:30]
        pageTableReg_1_0 <= io_cpu_din[4:0]; // @[NMK112.scala 91:30]
      end
    end
    if (io_cpu_wr) begin // @[NMK112.scala 88:19]
      if (chip & 2'h1 == bank) begin // @[NMK112.scala 91:30]
        pageTableReg_1_1 <= io_cpu_din[4:0]; // @[NMK112.scala 91:30]
      end
    end
    if (io_cpu_wr) begin // @[NMK112.scala 88:19]
      if (chip & 2'h2 == bank) begin // @[NMK112.scala 91:30]
        pageTableReg_1_2 <= io_cpu_din[4:0]; // @[NMK112.scala 91:30]
      end
    end
    if (io_cpu_wr) begin // @[NMK112.scala 88:19]
      if (chip & 2'h3 == bank) begin // @[NMK112.scala 91:30]
        pageTableReg_1_3 <= io_cpu_din[4:0]; // @[NMK112.scala 91:30]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pageTableReg_0_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  pageTableReg_0_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  pageTableReg_0_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  pageTableReg_0_3 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  pageTableReg_1_0 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  pageTableReg_1_1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  pageTableReg_1_2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  pageTableReg_1_3 = _RAND_7[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module OKIM6295(
  input         clock,
  input         reset,
  input         io_cpu_wr,
  input  [7:0]  io_cpu_din,
  output [7:0]  io_cpu_dout,
  output [17:0] io_rom_addr,
  input  [7:0]  io_rom_dout,
  input         io_rom_valid,
  output        io_audio_valid,
  output [13:0] io_audio_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  adpcm_rst; // @[OKIM6295.scala 96:21]
  wire  adpcm_clk; // @[OKIM6295.scala 96:21]
  wire  adpcm_cen; // @[OKIM6295.scala 96:21]
  wire  adpcm_ss; // @[OKIM6295.scala 96:21]
  wire  adpcm_wrn; // @[OKIM6295.scala 96:21]
  wire [7:0] adpcm_din; // @[OKIM6295.scala 96:21]
  wire [7:0] adpcm_dout; // @[OKIM6295.scala 96:21]
  wire [17:0] adpcm_rom_addr; // @[OKIM6295.scala 96:21]
  wire [7:0] adpcm_rom_data; // @[OKIM6295.scala 96:21]
  wire  adpcm_rom_ok; // @[OKIM6295.scala 96:21]
  wire [13:0] adpcm_sound; // @[OKIM6295.scala 96:21]
  wire  adpcm_sample; // @[OKIM6295.scala 96:21]
  reg [15:0] adpcm_io_cen_counter; // @[ClockDivider.scala 40:24]
  wire [16:0] adpcm_io_cen_next = adpcm_io_cen_counter + 16'h873; // @[ClockDivider.scala 42:19]
  reg  adpcm_io_cen_clockEnable; // @[ClockDivider.scala 41:28]
  jt6295 adpcm ( // @[OKIM6295.scala 96:21]
    .rst(adpcm_rst),
    .clk(adpcm_clk),
    .cen(adpcm_cen),
    .ss(adpcm_ss),
    .wrn(adpcm_wrn),
    .din(adpcm_din),
    .dout(adpcm_dout),
    .rom_addr(adpcm_rom_addr),
    .rom_data(adpcm_rom_data),
    .rom_ok(adpcm_rom_ok),
    .sound(adpcm_sound),
    .sample(adpcm_sample)
  );
  assign io_cpu_dout = adpcm_dout; // @[OKIM6295.scala 104:15]
  assign io_rom_addr = adpcm_rom_addr; // @[OKIM6295.scala 107:15]
  assign io_audio_valid = adpcm_sample; // @[OKIM6295.scala 111:18]
  assign io_audio_bits = adpcm_sound; // @[OKIM6295.scala 112:17]
  assign adpcm_rst = reset; // @[OKIM6295.scala 97:25]
  assign adpcm_clk = clock; // @[OKIM6295.scala 98:25]
  assign adpcm_cen = adpcm_io_cen_clockEnable; // @[OKIM6295.scala 99:16]
  assign adpcm_ss = 1'h1; // @[OKIM6295.scala 100:15]
  assign adpcm_wrn = ~io_cpu_wr; // @[OKIM6295.scala 102:19]
  assign adpcm_din = io_cpu_din; // @[OKIM6295.scala 103:16]
  assign adpcm_rom_data = io_rom_dout; // @[OKIM6295.scala 108:21]
  assign adpcm_rom_ok = io_rom_valid; // @[OKIM6295.scala 109:19]
  always @(posedge clock) begin
    adpcm_io_cen_counter <= adpcm_io_cen_counter + 16'h873; // @[ClockDivider.scala 40:34]
    adpcm_io_cen_clockEnable <= adpcm_io_cen_next[16]; // @[ClockDivider.scala 41:38]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  adpcm_io_cen_counter = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  adpcm_io_cen_clockEnable = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module OKIM6295_1(
  input         clock,
  input         reset,
  input         io_cpu_wr,
  input  [7:0]  io_cpu_din,
  output [7:0]  io_cpu_dout,
  output [17:0] io_rom_addr,
  input  [7:0]  io_rom_dout,
  input         io_rom_valid,
  output        io_audio_valid,
  output [13:0] io_audio_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  adpcm_rst; // @[OKIM6295.scala 96:21]
  wire  adpcm_clk; // @[OKIM6295.scala 96:21]
  wire  adpcm_cen; // @[OKIM6295.scala 96:21]
  wire  adpcm_ss; // @[OKIM6295.scala 96:21]
  wire  adpcm_wrn; // @[OKIM6295.scala 96:21]
  wire [7:0] adpcm_din; // @[OKIM6295.scala 96:21]
  wire [7:0] adpcm_dout; // @[OKIM6295.scala 96:21]
  wire [17:0] adpcm_rom_addr; // @[OKIM6295.scala 96:21]
  wire [7:0] adpcm_rom_data; // @[OKIM6295.scala 96:21]
  wire  adpcm_rom_ok; // @[OKIM6295.scala 96:21]
  wire [13:0] adpcm_sound; // @[OKIM6295.scala 96:21]
  wire  adpcm_sample; // @[OKIM6295.scala 96:21]
  reg [15:0] adpcm_io_cen_counter; // @[ClockDivider.scala 40:24]
  wire [16:0] adpcm_io_cen_next = adpcm_io_cen_counter + 16'h10e5; // @[ClockDivider.scala 42:19]
  reg  adpcm_io_cen_clockEnable; // @[ClockDivider.scala 41:28]
  jt6295 adpcm ( // @[OKIM6295.scala 96:21]
    .rst(adpcm_rst),
    .clk(adpcm_clk),
    .cen(adpcm_cen),
    .ss(adpcm_ss),
    .wrn(adpcm_wrn),
    .din(adpcm_din),
    .dout(adpcm_dout),
    .rom_addr(adpcm_rom_addr),
    .rom_data(adpcm_rom_data),
    .rom_ok(adpcm_rom_ok),
    .sound(adpcm_sound),
    .sample(adpcm_sample)
  );
  assign io_cpu_dout = adpcm_dout; // @[OKIM6295.scala 104:15]
  assign io_rom_addr = adpcm_rom_addr; // @[OKIM6295.scala 107:15]
  assign io_audio_valid = adpcm_sample; // @[OKIM6295.scala 111:18]
  assign io_audio_bits = adpcm_sound; // @[OKIM6295.scala 112:17]
  assign adpcm_rst = reset; // @[OKIM6295.scala 97:25]
  assign adpcm_clk = clock; // @[OKIM6295.scala 98:25]
  assign adpcm_cen = adpcm_io_cen_clockEnable; // @[OKIM6295.scala 99:16]
  assign adpcm_ss = 1'h1; // @[OKIM6295.scala 100:15]
  assign adpcm_wrn = ~io_cpu_wr; // @[OKIM6295.scala 102:19]
  assign adpcm_din = io_cpu_din; // @[OKIM6295.scala 103:16]
  assign adpcm_rom_data = io_rom_dout; // @[OKIM6295.scala 108:21]
  assign adpcm_rom_ok = io_rom_valid; // @[OKIM6295.scala 109:19]
  always @(posedge clock) begin
    adpcm_io_cen_counter <= adpcm_io_cen_counter + 16'h10e5; // @[ClockDivider.scala 40:34]
    adpcm_io_cen_clockEnable <= adpcm_io_cen_next[16]; // @[ClockDivider.scala 41:38]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  adpcm_io_cen_counter = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  adpcm_io_cen_clockEnable = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ADPCM(
  input  [3:0]  io_data,
  input  [16:0] io_in_step,
  input  [16:0] io_in_sample,
  output [16:0] io_out_step,
  output [16:0] io_out_sample
);
  wire [10:0] _GEN_4 = 3'h4 == io_data[2:0] ? $signed(11'sh133) : $signed(11'she6); // @[ADPCM.scala 75:{27,27}]
  wire [10:0] _GEN_5 = 3'h5 == io_data[2:0] ? $signed(11'sh199) : $signed(_GEN_4); // @[ADPCM.scala 75:{27,27}]
  wire [10:0] _GEN_6 = 3'h6 == io_data[2:0] ? $signed(11'sh200) : $signed(_GEN_5); // @[ADPCM.scala 75:{27,27}]
  wire [10:0] _GEN_7 = 3'h7 == io_data[2:0] ? $signed(11'sh266) : $signed(_GEN_6); // @[ADPCM.scala 75:{27,27}]
  wire [27:0] _step_T_1 = $signed(io_in_step) * $signed(_GEN_7); // @[ADPCM.scala 75:27]
  wire [19:0] step = _step_T_1[27:8]; // @[ADPCM.scala 75:48]
  wire [19:0] _io_out_step_T_1 = $signed(step) < 20'sh7f ? $signed(20'sh7f) : $signed(step); // @[Util.scala 264:51]
  wire [19:0] _io_out_step_T_3 = $signed(_io_out_step_T_1) < 20'sh6000 ? $signed(_io_out_step_T_1) : $signed(20'sh6000); // @[Util.scala 264:60]
  wire [4:0] _GEN_9 = 4'h1 == io_data ? $signed(5'sh3) : $signed(5'sh1); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_10 = 4'h2 == io_data ? $signed(5'sh5) : $signed(_GEN_9); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_11 = 4'h3 == io_data ? $signed(5'sh7) : $signed(_GEN_10); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_12 = 4'h4 == io_data ? $signed(5'sh9) : $signed(_GEN_11); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_13 = 4'h5 == io_data ? $signed(5'shb) : $signed(_GEN_12); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_14 = 4'h6 == io_data ? $signed(5'shd) : $signed(_GEN_13); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_15 = 4'h7 == io_data ? $signed(5'shf) : $signed(_GEN_14); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_16 = 4'h8 == io_data ? $signed(-5'sh1) : $signed(_GEN_15); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_17 = 4'h9 == io_data ? $signed(-5'sh3) : $signed(_GEN_16); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_18 = 4'ha == io_data ? $signed(-5'sh5) : $signed(_GEN_17); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_19 = 4'hb == io_data ? $signed(-5'sh7) : $signed(_GEN_18); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_20 = 4'hc == io_data ? $signed(-5'sh9) : $signed(_GEN_19); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_21 = 4'hd == io_data ? $signed(-5'shb) : $signed(_GEN_20); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_22 = 4'he == io_data ? $signed(-5'shd) : $signed(_GEN_21); // @[ADPCM.scala 79:{28,28}]
  wire [4:0] _GEN_23 = 4'hf == io_data ? $signed(-5'shf) : $signed(_GEN_22); // @[ADPCM.scala 79:{28,28}]
  wire [21:0] _delta_T = $signed(io_in_step) * $signed(_GEN_23); // @[ADPCM.scala 79:28]
  wire [18:0] delta = _delta_T[21:3]; // @[ADPCM.scala 79:50]
  wire [18:0] _GEN_24 = {{2{io_in_sample[16]}},io_in_sample}; // @[ADPCM.scala 80:44]
  wire [19:0] _io_out_sample_T = $signed(_GEN_24) + $signed(delta); // @[ADPCM.scala 80:44]
  wire [19:0] _io_out_sample_T_2 = $signed(_io_out_sample_T) < -20'sh8000 ? $signed(-20'sh8000) : $signed(
    _io_out_sample_T); // @[Util.scala 264:51]
  wire [19:0] _io_out_sample_T_4 = $signed(_io_out_sample_T_2) < 20'sh7fff ? $signed(_io_out_sample_T_2) : $signed(20'sh7fff
    ); // @[Util.scala 264:60]
  assign io_out_step = _io_out_step_T_3[16:0]; // @[ADPCM.scala 76:15]
  assign io_out_sample = _io_out_sample_T_4[16:0]; // @[ADPCM.scala 80:17]
endmodule
module LERP(
  input  [16:0] io_samples_0,
  input  [16:0] io_samples_1,
  input  [9:0]  io_index,
  output [16:0] io_out
);
  wire [17:0] slope = $signed(io_samples_1) - $signed(io_samples_0); // @[LERP.scala 54:29]
  wire [10:0] _offset_T = {1'b0,$signed(io_index)}; // @[LERP.scala 55:25]
  wire [28:0] _offset_T_1 = $signed(slope) * $signed(_offset_T); // @[LERP.scala 55:25]
  wire [27:0] offset = _offset_T_1[27:0]; // @[LERP.scala 55:25]
  wire [16:0] _io_out_T_1 = offset[25:9]; // @[LERP.scala 56:66]
  assign io_out = $signed(_io_out_T_1) + $signed(io_samples_0); // @[LERP.scala 56:73]
endmodule
module AudioPipeline(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits_state_samples_0,
  input  [15:0] io_in_bits_state_samples_1,
  input         io_in_bits_state_underflow,
  input  [15:0] io_in_bits_state_adpcmStep,
  input  [9:0]  io_in_bits_state_lerpIndex,
  input         io_in_bits_state_loopEnable,
  input  [15:0] io_in_bits_state_loopStep,
  input  [15:0] io_in_bits_state_loopSample,
  input  [7:0]  io_in_bits_pitch,
  input  [7:0]  io_in_bits_level,
  input  [3:0]  io_in_bits_pan,
  output        io_out_valid,
  output [15:0] io_out_bits_state_samples_0,
  output [15:0] io_out_bits_state_samples_1,
  output        io_out_bits_state_underflow,
  output [15:0] io_out_bits_state_adpcmStep,
  output [9:0]  io_out_bits_state_lerpIndex,
  output        io_out_bits_state_loopEnable,
  output [15:0] io_out_bits_state_loopStep,
  output [15:0] io_out_bits_state_loopSample,
  output [16:0] io_out_bits_audio_left,
  output        io_pcmData_ready,
  input         io_pcmData_valid,
  input  [3:0]  io_pcmData_bits,
  input         io_loopStart
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] adpcm_io_data; // @[AudioPipeline.scala 104:21]
  wire [16:0] adpcm_io_in_step; // @[AudioPipeline.scala 104:21]
  wire [16:0] adpcm_io_in_sample; // @[AudioPipeline.scala 104:21]
  wire [16:0] adpcm_io_out_step; // @[AudioPipeline.scala 104:21]
  wire [16:0] adpcm_io_out_sample; // @[AudioPipeline.scala 104:21]
  wire [16:0] lerp_io_samples_0; // @[AudioPipeline.scala 113:20]
  wire [16:0] lerp_io_samples_1; // @[AudioPipeline.scala 113:20]
  wire [9:0] lerp_io_index; // @[AudioPipeline.scala 113:20]
  wire [16:0] lerp_io_out; // @[AudioPipeline.scala 113:20]
  reg [2:0] stateReg; // @[AudioPipeline.scala 97:25]
  wire  _inputReg_T = io_in_ready & io_in_valid; // @[Decoupled.scala 52:35]
  reg [15:0] inputReg_state_samples_0; // @[Reg.scala 19:16]
  reg [15:0] inputReg_state_samples_1; // @[Reg.scala 19:16]
  reg  inputReg_state_underflow; // @[Reg.scala 19:16]
  reg [15:0] inputReg_state_adpcmStep; // @[Reg.scala 19:16]
  reg [9:0] inputReg_state_lerpIndex; // @[Reg.scala 19:16]
  reg  inputReg_state_loopEnable; // @[Reg.scala 19:16]
  reg [15:0] inputReg_state_loopStep; // @[Reg.scala 19:16]
  reg [15:0] inputReg_state_loopSample; // @[Reg.scala 19:16]
  reg [7:0] inputReg_pitch; // @[Reg.scala 19:16]
  reg [7:0] inputReg_level; // @[Reg.scala 19:16]
  reg [3:0] inputReg_pan; // @[Reg.scala 19:16]
  wire [15:0] _GEN_0 = _inputReg_T ? $signed(io_in_bits_state_samples_0) : $signed(inputReg_state_samples_0); // @[Reg.scala 19:16 20:{18,22}]
  wire [15:0] _GEN_1 = _inputReg_T ? $signed(io_in_bits_state_samples_1) : $signed(inputReg_state_samples_1); // @[Reg.scala 19:16 20:{18,22}]
  wire [15:0] _GEN_3 = _inputReg_T ? $signed(io_in_bits_state_adpcmStep) : $signed(inputReg_state_adpcmStep); // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_5 = _inputReg_T ? io_in_bits_state_loopEnable : inputReg_state_loopEnable; // @[Reg.scala 19:16 20:{18,22}]
  wire [15:0] _GEN_6 = _inputReg_T ? $signed(io_in_bits_state_loopStep) : $signed(inputReg_state_loopStep); // @[Reg.scala 19:16 20:{18,22}]
  wire [15:0] _GEN_7 = _inputReg_T ? $signed(io_in_bits_state_loopSample) : $signed(inputReg_state_loopSample); // @[Reg.scala 19:16 20:{18,22}]
  reg [16:0] sampleReg; // @[AudioPipeline.scala 99:22]
  reg [16:0] audioReg_left; // @[AudioPipeline.scala 100:21]
  wire  _pcmDataReg_T = io_pcmData_ready & io_pcmData_valid; // @[Decoupled.scala 52:35]
  reg [3:0] pcmDataReg; // @[Reg.scala 19:16]
  wire  _GEN_12 = io_loopStart & ~inputReg_state_loopEnable | _GEN_5; // @[AudioPipeline.scala 126:54 127:33]
  wire [16:0] _GEN_13 = io_loopStart & ~inputReg_state_loopEnable ? $signed(adpcm_io_out_step) : $signed({{1{_GEN_6[15
    ]}},_GEN_6}); // @[AudioPipeline.scala 126:54 128:31]
  wire [16:0] _GEN_14 = io_loopStart & ~inputReg_state_loopEnable ? $signed(adpcm_io_out_sample) : $signed({{1{_GEN_7[15
    ]}},_GEN_7}); // @[AudioPipeline.scala 126:54 129:33]
  wire  _step_T = io_loopStart & inputReg_state_loopEnable; // @[AudioPipeline.scala 131:33]
  wire [16:0] step = io_loopStart & inputReg_state_loopEnable ? $signed({{1{inputReg_state_loopStep[15]}},
    inputReg_state_loopStep}) : $signed(adpcm_io_out_step); // @[AudioPipeline.scala 131:19]
  wire [16:0] sample = _step_T ? $signed({{1{inputReg_state_loopSample[15]}},inputReg_state_loopSample}) : $signed(
    adpcm_io_out_sample); // @[AudioPipeline.scala 132:21]
  wire [16:0] _GEN_16 = stateReg == 3'h3 ? $signed(_GEN_13) : $signed({{1{_GEN_6[15]}},_GEN_6}); // @[AudioPipeline.scala 125:35]
  wire [16:0] _GEN_17 = stateReg == 3'h3 ? $signed(_GEN_14) : $signed({{1{_GEN_7[15]}},_GEN_7}); // @[AudioPipeline.scala 125:35]
  wire [16:0] _GEN_18 = stateReg == 3'h3 ? $signed(step) : $signed({{1{_GEN_3[15]}},_GEN_3}); // @[AudioPipeline.scala 125:35 AudioPipelineState.scala 57:15]
  wire [16:0] _WIRE_0 = {{1{inputReg_state_samples_1[15]}},inputReg_state_samples_1}; // @[AudioPipelineState.scala 58:{23,23}]
  wire [16:0] _GEN_19 = stateReg == 3'h3 ? $signed(_WIRE_0) : $signed({{1{_GEN_0[15]}},_GEN_0}); // @[AudioPipeline.scala 125:35 AudioPipelineState.scala 58:13]
  wire [16:0] _GEN_20 = stateReg == 3'h3 ? $signed(sample) : $signed({{1{_GEN_1[15]}},_GEN_1}); // @[AudioPipeline.scala 125:35 AudioPipelineState.scala 58:13]
  wire [9:0] _GEN_40 = {{2'd0}, inputReg_pitch}; // @[AudioPipelineState.scala 63:27]
  wire [9:0] _index_T_1 = inputReg_state_lerpIndex + _GEN_40; // @[AudioPipelineState.scala 63:27]
  wire [9:0] index = _index_T_1 + 10'h1; // @[AudioPipelineState.scala 63:35]
  wire [8:0] _sampleReg_T = inputReg_level + 8'h1; // @[AudioPipeline.scala 144:46]
  wire [9:0] _sampleReg_T_1 = {1'b0,$signed(_sampleReg_T)}; // @[AudioPipeline.scala 144:28]
  wire [26:0] _sampleReg_T_2 = $signed(sampleReg) * $signed(_sampleReg_T_1); // @[AudioPipeline.scala 144:28]
  wire [25:0] _sampleReg_T_4 = _sampleReg_T_2[25:0]; // @[AudioPipeline.scala 144:28]
  wire [16:0] _sampleReg_T_5 = _sampleReg_T_4[25:9]; // @[AudioPipeline.scala 144:54]
  wire [2:0] t = inputReg_pan[2:0]; // @[AudioPipeline.scala 150:25]
  wire [2:0] _left_T = ~t; // @[AudioPipeline.scala 156:20]
  wire [3:0] _left_T_1 = {1'b0,$signed(_left_T)}; // @[AudioPipeline.scala 156:17]
  wire [20:0] _left_T_2 = $signed(sampleReg) * $signed(_left_T_1); // @[AudioPipeline.scala 156:17]
  wire [19:0] _left_T_4 = _left_T_2[19:0]; // @[AudioPipeline.scala 156:17]
  wire [16:0] _left_T_5 = _left_T_4[19:3]; // @[AudioPipeline.scala 156:31]
  wire [2:0] _GEN_31 = io_pcmData_valid ? 3'h3 : stateReg; // @[AudioPipeline.scala 175:{30,41} 97:25]
  wire [2:0] _GEN_32 = 3'h7 == stateReg ? 3'h0 : stateReg; // @[AudioPipeline.scala 164:20 191:31 97:25]
  wire [2:0] _GEN_33 = 3'h6 == stateReg ? 3'h7 : _GEN_32; // @[AudioPipeline.scala 164:20 188:30]
  wire [2:0] _GEN_34 = 3'h5 == stateReg ? 3'h6 : _GEN_33; // @[AudioPipeline.scala 164:20 185:32]
  wire [2:0] _GEN_35 = 3'h4 == stateReg ? 3'h5 : _GEN_34; // @[AudioPipeline.scala 164:20 182:38]
  wire [2:0] _GEN_36 = 3'h3 == stateReg ? 3'h4 : _GEN_35; // @[AudioPipeline.scala 164:20 179:33]
  ADPCM adpcm ( // @[AudioPipeline.scala 104:21]
    .io_data(adpcm_io_data),
    .io_in_step(adpcm_io_in_step),
    .io_in_sample(adpcm_io_in_sample),
    .io_out_step(adpcm_io_out_step),
    .io_out_sample(adpcm_io_out_sample)
  );
  LERP lerp ( // @[AudioPipeline.scala 113:20]
    .io_samples_0(lerp_io_samples_0),
    .io_samples_1(lerp_io_samples_1),
    .io_index(lerp_io_index),
    .io_out(lerp_io_out)
  );
  assign io_in_ready = stateReg == 3'h0; // @[AudioPipeline.scala 195:27]
  assign io_out_valid = stateReg == 3'h7; // @[AudioPipeline.scala 196:28]
  assign io_out_bits_state_samples_0 = inputReg_state_samples_0; // @[AudioPipeline.scala 197:21]
  assign io_out_bits_state_samples_1 = inputReg_state_samples_1; // @[AudioPipeline.scala 197:21]
  assign io_out_bits_state_underflow = inputReg_state_underflow; // @[AudioPipeline.scala 197:21]
  assign io_out_bits_state_adpcmStep = inputReg_state_adpcmStep; // @[AudioPipeline.scala 197:21]
  assign io_out_bits_state_lerpIndex = inputReg_state_lerpIndex; // @[AudioPipeline.scala 197:21]
  assign io_out_bits_state_loopEnable = inputReg_state_loopEnable; // @[AudioPipeline.scala 197:21]
  assign io_out_bits_state_loopStep = inputReg_state_loopStep; // @[AudioPipeline.scala 197:21]
  assign io_out_bits_state_loopSample = inputReg_state_loopSample; // @[AudioPipeline.scala 197:21]
  assign io_out_bits_audio_left = audioReg_left; // @[AudioPipeline.scala 198:21]
  assign io_pcmData_ready = stateReg == 3'h2; // @[AudioPipeline.scala 199:32]
  assign adpcm_io_data = pcmDataReg; // @[AudioPipeline.scala 108:17]
  assign adpcm_io_in_step = {{1{inputReg_state_adpcmStep[15]}},inputReg_state_adpcmStep}; // @[AudioPipeline.scala 109:20]
  assign adpcm_io_in_sample = {{1{inputReg_state_samples_1[15]}},inputReg_state_samples_1}; // @[AudioPipeline.scala 110:22]
  assign lerp_io_samples_0 = {{1{inputReg_state_samples_0[15]}},inputReg_state_samples_0}; // @[AudioPipeline.scala 117:19]
  assign lerp_io_samples_1 = {{1{inputReg_state_samples_1[15]}},inputReg_state_samples_1}; // @[AudioPipeline.scala 117:19]
  assign lerp_io_index = inputReg_state_lerpIndex; // @[AudioPipeline.scala 118:17]
  always @(posedge clock) begin
    if (reset) begin // @[AudioPipeline.scala 97:25]
      stateReg <= 3'h0; // @[AudioPipeline.scala 97:25]
    end else if (3'h0 == stateReg) begin // @[AudioPipeline.scala 164:20]
      if (io_in_valid) begin // @[AudioPipeline.scala 167:25]
        stateReg <= 3'h1; // @[AudioPipeline.scala 167:36]
      end
    end else if (3'h1 == stateReg) begin // @[AudioPipeline.scala 164:20]
      if (inputReg_state_underflow) begin // @[AudioPipeline.scala 171:38]
        stateReg <= 3'h2;
      end else begin
        stateReg <= 3'h4;
      end
    end else if (3'h2 == stateReg) begin // @[AudioPipeline.scala 164:20]
      stateReg <= _GEN_31;
    end else begin
      stateReg <= _GEN_36;
    end
    inputReg_state_samples_0 <= _GEN_19[15:0];
    inputReg_state_samples_1 <= _GEN_20[15:0];
    if (stateReg == 3'h4) begin // @[AudioPipeline.scala 137:40]
      inputReg_state_underflow <= index[9]; // @[AudioPipelineState.scala 64:15]
    end else if (_inputReg_T) begin // @[Reg.scala 20:18]
      inputReg_state_underflow <= io_in_bits_state_underflow; // @[Reg.scala 20:22]
    end
    inputReg_state_adpcmStep <= _GEN_18[15:0];
    if (stateReg == 3'h4) begin // @[AudioPipeline.scala 137:40]
      inputReg_state_lerpIndex <= {{1'd0}, index[8:0]}; // @[AudioPipelineState.scala 65:15]
    end else if (_inputReg_T) begin // @[Reg.scala 20:18]
      inputReg_state_lerpIndex <= io_in_bits_state_lerpIndex; // @[Reg.scala 20:22]
    end
    if (stateReg == 3'h3) begin // @[AudioPipeline.scala 125:35]
      inputReg_state_loopEnable <= _GEN_12;
    end else if (_inputReg_T) begin // @[Reg.scala 20:18]
      inputReg_state_loopEnable <= io_in_bits_state_loopEnable; // @[Reg.scala 20:22]
    end
    inputReg_state_loopStep <= _GEN_16[15:0];
    inputReg_state_loopSample <= _GEN_17[15:0];
    if (_inputReg_T) begin // @[Reg.scala 20:18]
      inputReg_pitch <= io_in_bits_pitch; // @[Reg.scala 20:22]
    end
    if (_inputReg_T) begin // @[Reg.scala 20:18]
      inputReg_level <= io_in_bits_level; // @[Reg.scala 20:22]
    end
    if (_inputReg_T) begin // @[Reg.scala 20:18]
      inputReg_pan <= io_in_bits_pan; // @[Reg.scala 20:22]
    end
    if (stateReg == 3'h5) begin // @[AudioPipeline.scala 143:34]
      sampleReg <= _sampleReg_T_5; // @[AudioPipeline.scala 144:15]
    end else if (stateReg == 3'h4) begin // @[AudioPipeline.scala 137:40]
      sampleReg <= lerp_io_out; // @[AudioPipeline.scala 139:15]
    end
    if (stateReg == 3'h6) begin // @[AudioPipeline.scala 148:32]
      if (inputReg_pan > 4'h8) begin // @[AudioPipeline.scala 155:30]
        audioReg_left <= _left_T_5; // @[AudioPipeline.scala 156:12]
      end else begin
        audioReg_left <= sampleReg; // @[AudioPipeline.scala 153:10]
      end
    end
    if (_pcmDataReg_T) begin // @[Reg.scala 20:18]
      pcmDataReg <= io_pcmData_bits; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  inputReg_state_samples_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  inputReg_state_samples_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  inputReg_state_underflow = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  inputReg_state_adpcmStep = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  inputReg_state_lerpIndex = _RAND_5[9:0];
  _RAND_6 = {1{`RANDOM}};
  inputReg_state_loopEnable = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  inputReg_state_loopStep = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  inputReg_state_loopSample = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  inputReg_pitch = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  inputReg_level = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  inputReg_pan = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  sampleReg = _RAND_12[16:0];
  _RAND_13 = {1{`RANDOM}};
  audioReg_left = _RAND_13[16:0];
  _RAND_14 = {1{`RANDOM}};
  pcmDataReg = _RAND_14[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ChannelController(
  input         clock,
  input         reset,
  input  [7:0]  io_regs_0_pitch,
  input         io_regs_0_flags_keyOn,
  input         io_regs_0_flags_loop,
  input  [7:0]  io_regs_0_level,
  input  [3:0]  io_regs_0_pan,
  input  [23:0] io_regs_0_startAddr,
  input  [23:0] io_regs_0_loopStartAddr,
  input  [23:0] io_regs_0_loopEndAddr,
  input  [23:0] io_regs_0_endAddr,
  input  [7:0]  io_regs_1_pitch,
  input         io_regs_1_flags_keyOn,
  input         io_regs_1_flags_loop,
  input  [7:0]  io_regs_1_level,
  input  [3:0]  io_regs_1_pan,
  input  [23:0] io_regs_1_startAddr,
  input  [23:0] io_regs_1_loopStartAddr,
  input  [23:0] io_regs_1_loopEndAddr,
  input  [23:0] io_regs_1_endAddr,
  input  [7:0]  io_regs_2_pitch,
  input         io_regs_2_flags_keyOn,
  input         io_regs_2_flags_loop,
  input  [7:0]  io_regs_2_level,
  input  [3:0]  io_regs_2_pan,
  input  [23:0] io_regs_2_startAddr,
  input  [23:0] io_regs_2_loopStartAddr,
  input  [23:0] io_regs_2_loopEndAddr,
  input  [23:0] io_regs_2_endAddr,
  input  [7:0]  io_regs_3_pitch,
  input         io_regs_3_flags_keyOn,
  input         io_regs_3_flags_loop,
  input  [7:0]  io_regs_3_level,
  input  [3:0]  io_regs_3_pan,
  input  [23:0] io_regs_3_startAddr,
  input  [23:0] io_regs_3_loopStartAddr,
  input  [23:0] io_regs_3_loopEndAddr,
  input  [23:0] io_regs_3_endAddr,
  input  [7:0]  io_regs_4_pitch,
  input         io_regs_4_flags_keyOn,
  input         io_regs_4_flags_loop,
  input  [7:0]  io_regs_4_level,
  input  [3:0]  io_regs_4_pan,
  input  [23:0] io_regs_4_startAddr,
  input  [23:0] io_regs_4_loopStartAddr,
  input  [23:0] io_regs_4_loopEndAddr,
  input  [23:0] io_regs_4_endAddr,
  input  [7:0]  io_regs_5_pitch,
  input         io_regs_5_flags_keyOn,
  input         io_regs_5_flags_loop,
  input  [7:0]  io_regs_5_level,
  input  [3:0]  io_regs_5_pan,
  input  [23:0] io_regs_5_startAddr,
  input  [23:0] io_regs_5_loopStartAddr,
  input  [23:0] io_regs_5_loopEndAddr,
  input  [23:0] io_regs_5_endAddr,
  input  [7:0]  io_regs_6_pitch,
  input         io_regs_6_flags_keyOn,
  input         io_regs_6_flags_loop,
  input  [7:0]  io_regs_6_level,
  input  [3:0]  io_regs_6_pan,
  input  [23:0] io_regs_6_startAddr,
  input  [23:0] io_regs_6_loopStartAddr,
  input  [23:0] io_regs_6_loopEndAddr,
  input  [23:0] io_regs_6_endAddr,
  input  [7:0]  io_regs_7_pitch,
  input         io_regs_7_flags_keyOn,
  input         io_regs_7_flags_loop,
  input  [7:0]  io_regs_7_level,
  input  [3:0]  io_regs_7_pan,
  input  [23:0] io_regs_7_startAddr,
  input  [23:0] io_regs_7_loopStartAddr,
  input  [23:0] io_regs_7_loopEndAddr,
  input  [23:0] io_regs_7_endAddr,
  input         io_enable,
  output        io_done,
  output [2:0]  io_index,
  output        io_audio_valid,
  output [15:0] io_audio_bits_left,
  output        io_rom_rd,
  output [23:0] io_rom_addr,
  input  [7:0]  io_rom_dout,
  input         io_rom_wait_n,
  input         io_rom_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] channelStateMem [0:7]; // @[ChannelController.scala 99:36]
  wire  channelStateMem_channelState_MPORT_en; // @[ChannelController.scala 99:36]
  wire [2:0] channelStateMem_channelState_MPORT_addr; // @[ChannelController.scala 99:36]
  wire [120:0] channelStateMem_channelState_MPORT_data; // @[ChannelController.scala 99:36]
  wire [120:0] channelStateMem_MPORT_data; // @[ChannelController.scala 99:36]
  wire [2:0] channelStateMem_MPORT_addr; // @[ChannelController.scala 99:36]
  wire  channelStateMem_MPORT_mask; // @[ChannelController.scala 99:36]
  wire  channelStateMem_MPORT_en; // @[ChannelController.scala 99:36]
  reg  channelStateMem_channelState_MPORT_en_pipe_0;
  reg [2:0] channelStateMem_channelState_MPORT_addr_pipe_0;
  wire  audioPipeline_clock; // @[ChannelController.scala 104:29]
  wire  audioPipeline_reset; // @[ChannelController.scala 104:29]
  wire  audioPipeline_io_in_ready; // @[ChannelController.scala 104:29]
  wire  audioPipeline_io_in_valid; // @[ChannelController.scala 104:29]
  wire [15:0] audioPipeline_io_in_bits_state_samples_0; // @[ChannelController.scala 104:29]
  wire [15:0] audioPipeline_io_in_bits_state_samples_1; // @[ChannelController.scala 104:29]
  wire  audioPipeline_io_in_bits_state_underflow; // @[ChannelController.scala 104:29]
  wire [15:0] audioPipeline_io_in_bits_state_adpcmStep; // @[ChannelController.scala 104:29]
  wire [9:0] audioPipeline_io_in_bits_state_lerpIndex; // @[ChannelController.scala 104:29]
  wire  audioPipeline_io_in_bits_state_loopEnable; // @[ChannelController.scala 104:29]
  wire [15:0] audioPipeline_io_in_bits_state_loopStep; // @[ChannelController.scala 104:29]
  wire [15:0] audioPipeline_io_in_bits_state_loopSample; // @[ChannelController.scala 104:29]
  wire [7:0] audioPipeline_io_in_bits_pitch; // @[ChannelController.scala 104:29]
  wire [7:0] audioPipeline_io_in_bits_level; // @[ChannelController.scala 104:29]
  wire [3:0] audioPipeline_io_in_bits_pan; // @[ChannelController.scala 104:29]
  wire  audioPipeline_io_out_valid; // @[ChannelController.scala 104:29]
  wire [15:0] audioPipeline_io_out_bits_state_samples_0; // @[ChannelController.scala 104:29]
  wire [15:0] audioPipeline_io_out_bits_state_samples_1; // @[ChannelController.scala 104:29]
  wire  audioPipeline_io_out_bits_state_underflow; // @[ChannelController.scala 104:29]
  wire [15:0] audioPipeline_io_out_bits_state_adpcmStep; // @[ChannelController.scala 104:29]
  wire [9:0] audioPipeline_io_out_bits_state_lerpIndex; // @[ChannelController.scala 104:29]
  wire  audioPipeline_io_out_bits_state_loopEnable; // @[ChannelController.scala 104:29]
  wire [15:0] audioPipeline_io_out_bits_state_loopStep; // @[ChannelController.scala 104:29]
  wire [15:0] audioPipeline_io_out_bits_state_loopSample; // @[ChannelController.scala 104:29]
  wire [16:0] audioPipeline_io_out_bits_audio_left; // @[ChannelController.scala 104:29]
  wire  audioPipeline_io_pcmData_ready; // @[ChannelController.scala 104:29]
  wire  audioPipeline_io_pcmData_valid; // @[ChannelController.scala 104:29]
  wire [3:0] audioPipeline_io_pcmData_bits; // @[ChannelController.scala 104:29]
  wire  audioPipeline_io_loopStart; // @[ChannelController.scala 104:29]
  reg [3:0] stateReg; // @[ChannelController.scala 88:25]
  reg [16:0] accumulatorReg_left; // @[ChannelController.scala 89:27]
  wire  _T = stateReg == 4'h0; // @[ChannelController.scala 92:99]
  wire  _T_2 = stateReg == 4'h0 | stateReg == 4'h8; // @[ChannelController.scala 92:114]
  reg [2:0] channelCounter; // @[Counter.scala 40:34]
  wire  wrap_wrap = channelCounter == 3'h7; // @[Counter.scala 45:24]
  wire [2:0] _wrap_value_T_1 = channelCounter + 3'h1; // @[Counter.scala 46:22]
  wire  channelCounterWrap = _T_2 & wrap_wrap; // @[Counter.scala 86:{48,55}]
  reg [8:0] outputCounterWrap_value; // @[Counter.scala 40:34]
  wire  outputCounterWrap_wrap_wrap = outputCounterWrap_value == 9'h16a; // @[Counter.scala 45:24]
  wire [8:0] _outputCounterWrap_wrap_value_T_1 = outputCounterWrap_value + 9'h1; // @[Counter.scala 46:22]
  wire [120:0] _channelState_WIRE_1 = channelStateMem_channelState_MPORT_data;
  wire [15:0] channelState_audioPipelineState_loopSample = _channelState_WIRE_1[15:0]; // @[ChannelController.scala 100:92]
  wire [15:0] channelState_audioPipelineState_loopStep = _channelState_WIRE_1[31:16]; // @[ChannelController.scala 100:92]
  wire  channelState_audioPipelineState_loopEnable = _channelState_WIRE_1[32]; // @[ChannelController.scala 100:92]
  wire [9:0] channelState_audioPipelineState_lerpIndex = _channelState_WIRE_1[42:33]; // @[ChannelController.scala 100:92]
  wire [15:0] channelState_audioPipelineState_adpcmStep = _channelState_WIRE_1[58:43]; // @[ChannelController.scala 100:92]
  wire  channelState_audioPipelineState_underflow = _channelState_WIRE_1[59]; // @[ChannelController.scala 100:92]
  wire [15:0] channelState_audioPipelineState_samples_0 = _channelState_WIRE_1[75:60]; // @[ChannelController.scala 100:92]
  wire [15:0] channelState_audioPipelineState_samples_1 = _channelState_WIRE_1[91:76]; // @[ChannelController.scala 100:92]
  wire  channelState_loopStart = _channelState_WIRE_1[92]; // @[ChannelController.scala 100:92]
  wire [23:0] channelState_addr = _channelState_WIRE_1[116:93]; // @[ChannelController.scala 100:92]
  wire  channelState_nibble = _channelState_WIRE_1[117]; // @[ChannelController.scala 100:92]
  wire  channelState_done = _channelState_WIRE_1[118]; // @[ChannelController.scala 100:92]
  wire  channelState_active = _channelState_WIRE_1[119]; // @[ChannelController.scala 100:92]
  wire  channelState_enable = _channelState_WIRE_1[120]; // @[ChannelController.scala 100:92]
  wire  _channelStateReg_T = stateReg == 4'h3; // @[ChannelController.scala 101:58]
  reg  channelStateReg_enable; // @[Reg.scala 19:16]
  reg  channelStateReg_active; // @[Reg.scala 19:16]
  reg  channelStateReg_done; // @[Reg.scala 19:16]
  reg  channelStateReg_nibble; // @[Reg.scala 19:16]
  reg [23:0] channelStateReg_addr; // @[Reg.scala 19:16]
  reg  channelStateReg_loopStart; // @[Reg.scala 19:16]
  reg [15:0] channelStateReg_audioPipelineState_samples_0; // @[Reg.scala 19:16]
  reg [15:0] channelStateReg_audioPipelineState_samples_1; // @[Reg.scala 19:16]
  reg  channelStateReg_audioPipelineState_underflow; // @[Reg.scala 19:16]
  reg [15:0] channelStateReg_audioPipelineState_adpcmStep; // @[Reg.scala 19:16]
  reg [9:0] channelStateReg_audioPipelineState_lerpIndex; // @[Reg.scala 19:16]
  reg  channelStateReg_audioPipelineState_loopEnable; // @[Reg.scala 19:16]
  reg [15:0] channelStateReg_audioPipelineState_loopStep; // @[Reg.scala 19:16]
  reg [15:0] channelStateReg_audioPipelineState_loopSample; // @[Reg.scala 19:16]
  wire  _GEN_13 = _channelStateReg_T ? channelState_enable : channelStateReg_enable; // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_14 = _channelStateReg_T ? channelState_active : channelStateReg_active; // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_15 = _channelStateReg_T ? channelState_done : channelStateReg_done; // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_16 = _channelStateReg_T ? channelState_nibble : channelStateReg_nibble; // @[Reg.scala 19:16 20:{18,22}]
  wire [23:0] _GEN_17 = _channelStateReg_T ? channelState_addr : channelStateReg_addr; // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_18 = _channelStateReg_T ? channelState_loopStart : channelStateReg_loopStart; // @[Reg.scala 19:16 20:{18,22}]
  wire [15:0] _GEN_19 = _channelStateReg_T ? $signed(channelState_audioPipelineState_samples_0) : $signed(
    channelStateReg_audioPipelineState_samples_0); // @[Reg.scala 19:16 20:{18,22}]
  wire [15:0] _GEN_20 = _channelStateReg_T ? $signed(channelState_audioPipelineState_samples_1) : $signed(
    channelStateReg_audioPipelineState_samples_1); // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_21 = _channelStateReg_T ? channelState_audioPipelineState_underflow :
    channelStateReg_audioPipelineState_underflow; // @[Reg.scala 19:16 20:{18,22}]
  wire [15:0] _GEN_22 = _channelStateReg_T ? $signed(channelState_audioPipelineState_adpcmStep) : $signed(
    channelStateReg_audioPipelineState_adpcmStep); // @[Reg.scala 19:16 20:{18,22}]
  wire [9:0] _GEN_23 = _channelStateReg_T ? channelState_audioPipelineState_lerpIndex :
    channelStateReg_audioPipelineState_lerpIndex; // @[Reg.scala 19:16 20:{18,22}]
  wire  _GEN_24 = _channelStateReg_T ? channelState_audioPipelineState_loopEnable :
    channelStateReg_audioPipelineState_loopEnable; // @[Reg.scala 19:16 20:{18,22}]
  wire [15:0] _GEN_25 = _channelStateReg_T ? $signed(channelState_audioPipelineState_loopStep) : $signed(
    channelStateReg_audioPipelineState_loopStep); // @[Reg.scala 19:16 20:{18,22}]
  wire [15:0] _GEN_26 = _channelStateReg_T ? $signed(channelState_audioPipelineState_loopSample) : $signed(
    channelStateReg_audioPipelineState_loopSample); // @[Reg.scala 19:16 20:{18,22}]
  wire [7:0] _GEN_28 = 3'h1 == channelCounter ? io_regs_1_pitch : io_regs_0_pitch; // @[ChannelController.scala 107:{34,34}]
  wire [7:0] _GEN_29 = 3'h2 == channelCounter ? io_regs_2_pitch : _GEN_28; // @[ChannelController.scala 107:{34,34}]
  wire [7:0] _GEN_30 = 3'h3 == channelCounter ? io_regs_3_pitch : _GEN_29; // @[ChannelController.scala 107:{34,34}]
  wire [7:0] _GEN_31 = 3'h4 == channelCounter ? io_regs_4_pitch : _GEN_30; // @[ChannelController.scala 107:{34,34}]
  wire [7:0] _GEN_32 = 3'h5 == channelCounter ? io_regs_5_pitch : _GEN_31; // @[ChannelController.scala 107:{34,34}]
  wire [7:0] _GEN_33 = 3'h6 == channelCounter ? io_regs_6_pitch : _GEN_32; // @[ChannelController.scala 107:{34,34}]
  wire [7:0] _GEN_36 = 3'h1 == channelCounter ? io_regs_1_level : io_regs_0_level; // @[ChannelController.scala 108:{34,34}]
  wire [7:0] _GEN_37 = 3'h2 == channelCounter ? io_regs_2_level : _GEN_36; // @[ChannelController.scala 108:{34,34}]
  wire [7:0] _GEN_38 = 3'h3 == channelCounter ? io_regs_3_level : _GEN_37; // @[ChannelController.scala 108:{34,34}]
  wire [7:0] _GEN_39 = 3'h4 == channelCounter ? io_regs_4_level : _GEN_38; // @[ChannelController.scala 108:{34,34}]
  wire [7:0] _GEN_40 = 3'h5 == channelCounter ? io_regs_5_level : _GEN_39; // @[ChannelController.scala 108:{34,34}]
  wire [7:0] _GEN_41 = 3'h6 == channelCounter ? io_regs_6_level : _GEN_40; // @[ChannelController.scala 108:{34,34}]
  wire [3:0] _GEN_44 = 3'h1 == channelCounter ? io_regs_1_pan : io_regs_0_pan; // @[ChannelController.scala 109:{32,32}]
  wire [3:0] _GEN_45 = 3'h2 == channelCounter ? io_regs_2_pan : _GEN_44; // @[ChannelController.scala 109:{32,32}]
  wire [3:0] _GEN_46 = 3'h3 == channelCounter ? io_regs_3_pan : _GEN_45; // @[ChannelController.scala 109:{32,32}]
  wire [3:0] _GEN_47 = 3'h4 == channelCounter ? io_regs_4_pan : _GEN_46; // @[ChannelController.scala 109:{32,32}]
  wire [3:0] _GEN_48 = 3'h5 == channelCounter ? io_regs_5_pan : _GEN_47; // @[ChannelController.scala 109:{32,32}]
  wire [3:0] _GEN_49 = 3'h6 == channelCounter ? io_regs_6_pan : _GEN_48; // @[ChannelController.scala 109:{32,32}]
  wire  _GEN_52 = 3'h1 == channelCounter ? io_regs_1_flags_keyOn : io_regs_0_flags_keyOn; // @[ChannelController.scala 115:{66,66}]
  wire  _GEN_53 = 3'h2 == channelCounter ? io_regs_2_flags_keyOn : _GEN_52; // @[ChannelController.scala 115:{66,66}]
  wire  _GEN_54 = 3'h3 == channelCounter ? io_regs_3_flags_keyOn : _GEN_53; // @[ChannelController.scala 115:{66,66}]
  wire  _GEN_55 = 3'h4 == channelCounter ? io_regs_4_flags_keyOn : _GEN_54; // @[ChannelController.scala 115:{66,66}]
  wire  _GEN_56 = 3'h5 == channelCounter ? io_regs_5_flags_keyOn : _GEN_55; // @[ChannelController.scala 115:{66,66}]
  wire  _GEN_57 = 3'h6 == channelCounter ? io_regs_6_flags_keyOn : _GEN_56; // @[ChannelController.scala 115:{66,66}]
  wire  _GEN_58 = 3'h7 == channelCounter ? io_regs_7_flags_keyOn : _GEN_57; // @[ChannelController.scala 115:{66,66}]
  wire  start = ~channelStateReg_enable & ~channelStateReg_active & _GEN_58; // @[ChannelController.scala 115:66]
  wire  stop = channelStateReg_enable & ~_GEN_58; // @[ChannelController.scala 116:37]
  wire  active = channelStateReg_active | start; // @[ChannelController.scala 117:39]
  wire  _pendingReg_T = audioPipeline_io_pcmData_ready & io_rom_wait_n; // @[ChannelController.scala 121:66]
  reg  pendingReg; // @[Util.scala 218:28]
  wire  _GEN_59 = _pendingReg_T | pendingReg; // @[Util.scala 218:28 219:{54,66}]
  wire  _T_4 = stateReg == 4'h4; // @[ChannelController.scala 129:17]
  wire [23:0] _GEN_64 = 3'h1 == channelCounter ? io_regs_1_startAddr : io_regs_0_startAddr; // @[ChannelState.scala 61:{10,10}]
  wire [23:0] _GEN_65 = 3'h2 == channelCounter ? io_regs_2_startAddr : _GEN_64; // @[ChannelState.scala 61:{10,10}]
  wire [23:0] _GEN_66 = 3'h3 == channelCounter ? io_regs_3_startAddr : _GEN_65; // @[ChannelState.scala 61:{10,10}]
  wire [23:0] _GEN_67 = 3'h4 == channelCounter ? io_regs_4_startAddr : _GEN_66; // @[ChannelState.scala 61:{10,10}]
  wire [23:0] _GEN_68 = 3'h5 == channelCounter ? io_regs_5_startAddr : _GEN_67; // @[ChannelState.scala 61:{10,10}]
  wire [23:0] _GEN_69 = 3'h6 == channelCounter ? io_regs_6_startAddr : _GEN_68; // @[ChannelState.scala 61:{10,10}]
  wire [23:0] _GEN_70 = 3'h7 == channelCounter ? io_regs_7_startAddr : _GEN_69; // @[ChannelState.scala 61:{10,10}]
  wire  _GEN_71 = channelStateReg_done ? 1'h0 : _GEN_15; // @[ChannelController.scala 134:22 ChannelState.scala 97:10]
  wire  _GEN_72 = stop ? 1'h0 : _GEN_13; // @[ChannelController.scala 132:22 ChannelState.scala 68:12]
  wire  _GEN_73 = stop ? 1'h0 : _GEN_14; // @[ChannelController.scala 132:22 ChannelState.scala 69:12]
  wire  _GEN_74 = stop ? 1'h0 : _GEN_71; // @[ChannelController.scala 132:22 ChannelState.scala 70:10]
  wire  _GEN_75 = start | _GEN_72; // @[ChannelController.scala 130:17 ChannelState.scala 57:12]
  wire  _GEN_76 = start | _GEN_73; // @[ChannelController.scala 130:17 ChannelState.scala 58:12]
  wire  _GEN_77 = start ? 1'h0 : _GEN_74; // @[ChannelController.scala 130:17 ChannelState.scala 59:10]
  wire [23:0] _GEN_79 = start ? _GEN_70 : _GEN_17; // @[ChannelController.scala 130:17 ChannelState.scala 61:10]
  wire  _GEN_83 = start | _GEN_21; // @[ChannelController.scala 130:17 ChannelState.scala 63:24]
  wire  _GEN_90 = stateReg == 4'h4 ? _GEN_76 : _GEN_14; // @[ChannelController.scala 129:34]
  wire  _GEN_91 = stateReg == 4'h4 ? _GEN_77 : _GEN_15; // @[ChannelController.scala 129:34]
  wire [23:0] _GEN_93 = stateReg == 4'h4 ? _GEN_79 : _GEN_17; // @[ChannelController.scala 129:34]
  wire  _T_5 = audioPipeline_io_pcmData_ready & audioPipeline_io_pcmData_valid; // @[Decoupled.scala 52:35]
  wire [23:0] _GEN_104 = 3'h1 == channelCounter ? io_regs_1_loopStartAddr : io_regs_0_loopStartAddr; // @[ChannelState.scala 81:{48,48}]
  wire [23:0] _GEN_105 = 3'h2 == channelCounter ? io_regs_2_loopStartAddr : _GEN_104; // @[ChannelState.scala 81:{48,48}]
  wire [23:0] _GEN_106 = 3'h3 == channelCounter ? io_regs_3_loopStartAddr : _GEN_105; // @[ChannelState.scala 81:{48,48}]
  wire [23:0] _GEN_107 = 3'h4 == channelCounter ? io_regs_4_loopStartAddr : _GEN_106; // @[ChannelState.scala 81:{48,48}]
  wire [23:0] _GEN_108 = 3'h5 == channelCounter ? io_regs_5_loopStartAddr : _GEN_107; // @[ChannelState.scala 81:{48,48}]
  wire [23:0] _GEN_109 = 3'h6 == channelCounter ? io_regs_6_loopStartAddr : _GEN_108; // @[ChannelState.scala 81:{48,48}]
  wire [23:0] _GEN_110 = 3'h7 == channelCounter ? io_regs_7_loopStartAddr : _GEN_109; // @[ChannelState.scala 81:{48,48}]
  wire  _GEN_112 = 3'h1 == channelCounter ? io_regs_1_flags_loop : io_regs_0_flags_loop; // @[ChannelState.scala 81:{40,40}]
  wire  _GEN_113 = 3'h2 == channelCounter ? io_regs_2_flags_loop : _GEN_112; // @[ChannelState.scala 81:{40,40}]
  wire  _GEN_114 = 3'h3 == channelCounter ? io_regs_3_flags_loop : _GEN_113; // @[ChannelState.scala 81:{40,40}]
  wire  _GEN_115 = 3'h4 == channelCounter ? io_regs_4_flags_loop : _GEN_114; // @[ChannelState.scala 81:{40,40}]
  wire  _GEN_116 = 3'h5 == channelCounter ? io_regs_5_flags_loop : _GEN_115; // @[ChannelState.scala 81:{40,40}]
  wire  _GEN_117 = 3'h6 == channelCounter ? io_regs_6_flags_loop : _GEN_116; // @[ChannelState.scala 81:{40,40}]
  wire  _GEN_118 = 3'h7 == channelCounter ? io_regs_7_flags_loop : _GEN_117; // @[ChannelState.scala 81:{40,40}]
  wire  _channelStateReg_loopStart_T_2 = ~channelStateReg_nibble; // @[ChannelState.scala 81:80]
  wire [23:0] _GEN_120 = 3'h1 == channelCounter ? io_regs_1_loopEndAddr : io_regs_0_loopEndAddr; // @[ChannelState.scala 84:{42,42}]
  wire [23:0] _GEN_121 = 3'h2 == channelCounter ? io_regs_2_loopEndAddr : _GEN_120; // @[ChannelState.scala 84:{42,42}]
  wire [23:0] _GEN_122 = 3'h3 == channelCounter ? io_regs_3_loopEndAddr : _GEN_121; // @[ChannelState.scala 84:{42,42}]
  wire [23:0] _GEN_123 = 3'h4 == channelCounter ? io_regs_4_loopEndAddr : _GEN_122; // @[ChannelState.scala 84:{42,42}]
  wire [23:0] _GEN_124 = 3'h5 == channelCounter ? io_regs_5_loopEndAddr : _GEN_123; // @[ChannelState.scala 84:{42,42}]
  wire [23:0] _GEN_125 = 3'h6 == channelCounter ? io_regs_6_loopEndAddr : _GEN_124; // @[ChannelState.scala 84:{42,42}]
  wire [23:0] _GEN_126 = 3'h7 == channelCounter ? io_regs_7_loopEndAddr : _GEN_125; // @[ChannelState.scala 84:{42,42}]
  wire [23:0] _GEN_128 = 3'h1 == channelCounter ? io_regs_1_endAddr : io_regs_0_endAddr; // @[ChannelState.scala 86:{23,23}]
  wire [23:0] _GEN_129 = 3'h2 == channelCounter ? io_regs_2_endAddr : _GEN_128; // @[ChannelState.scala 86:{23,23}]
  wire [23:0] _GEN_130 = 3'h3 == channelCounter ? io_regs_3_endAddr : _GEN_129; // @[ChannelState.scala 86:{23,23}]
  wire [23:0] _GEN_131 = 3'h4 == channelCounter ? io_regs_4_endAddr : _GEN_130; // @[ChannelState.scala 86:{23,23}]
  wire [23:0] _GEN_132 = 3'h5 == channelCounter ? io_regs_5_endAddr : _GEN_131; // @[ChannelState.scala 86:{23,23}]
  wire [23:0] _GEN_133 = 3'h6 == channelCounter ? io_regs_6_endAddr : _GEN_132; // @[ChannelState.scala 86:{23,23}]
  wire [23:0] _GEN_134 = 3'h7 == channelCounter ? io_regs_7_endAddr : _GEN_133; // @[ChannelState.scala 86:{23,23}]
  wire [23:0] _channelStateReg_addr_T_1 = channelStateReg_addr + 24'h1; // @[ChannelState.scala 90:22]
  wire  _GEN_136 = channelStateReg_addr == _GEN_134 | _GEN_91; // @[ChannelState.scala 86:47 88:14]
  wire [16:0] accumulatorReg_sample_1_left = $signed(accumulatorReg_left) + $signed(audioPipeline_io_out_bits_audio_left
    ); // @[Audio.scala 51:47]
  wire  _T_10 = stateReg == 4'h7; // @[ChannelController.scala 152:44]
  wire  data_enable = _T_10 & channelStateReg_enable; // @[ChannelController.scala 153:19]
  wire  data_active = _T_10 & channelStateReg_active; // @[ChannelController.scala 153:19]
  wire  data_done = _T_10 & channelStateReg_done; // @[ChannelController.scala 153:19]
  wire  data_nibble = _T_10 & channelStateReg_nibble; // @[ChannelController.scala 153:19]
  wire [23:0] data_addr = _T_10 ? channelStateReg_addr : 24'h0; // @[ChannelController.scala 153:19]
  wire  data_loopStart = _T_10 & channelStateReg_loopStart; // @[ChannelController.scala 153:19]
  wire  data_audioPipelineState_underflow = _T_10 ? channelStateReg_audioPipelineState_underflow : 1'h1; // @[ChannelController.scala 153:19]
  wire [9:0] data_audioPipelineState_lerpIndex = _T_10 ? channelStateReg_audioPipelineState_lerpIndex : 10'h0; // @[ChannelController.scala 153:19]
  wire  data_audioPipelineState_loopEnable = _T_10 & channelStateReg_audioPipelineState_loopEnable; // @[ChannelController.scala 153:19]
  wire [15:0] _T_12 = _T_10 ? $signed(channelStateReg_audioPipelineState_loopSample) : $signed(16'sh0); // @[ChannelController.scala 154:48]
  wire [15:0] _T_13 = _T_10 ? $signed(channelStateReg_audioPipelineState_loopStep) : $signed(16'sh0); // @[ChannelController.scala 154:48]
  wire [15:0] _T_14 = _T_10 ? $signed(channelStateReg_audioPipelineState_adpcmStep) : $signed(16'sh7f); // @[ChannelController.scala 154:48]
  wire [15:0] _T_15 = _T_10 ? $signed(channelStateReg_audioPipelineState_samples_0) : $signed(16'sh0); // @[ChannelController.scala 154:48]
  wire [15:0] _T_16 = _T_10 ? $signed(channelStateReg_audioPipelineState_samples_1) : $signed(16'sh0); // @[ChannelController.scala 154:48]
  wire [75:0] lo = {_T_15,data_audioPipelineState_underflow,_T_14,data_audioPipelineState_lerpIndex,
    data_audioPipelineState_loopEnable,_T_13,_T_12}; // @[ChannelController.scala 154:48]
  wire [44:0] hi = {data_enable,data_active,data_done,data_nibble,data_addr,data_loopStart,_T_16}; // @[ChannelController.scala 154:48]
  wire [3:0] _stateReg_T = active ? 4'h5 : 4'h7; // @[ChannelController.scala 176:38]
  wire [3:0] _GEN_166 = audioPipeline_io_in_ready ? 4'h6 : stateReg; // @[ChannelController.scala 180:{39,50} 88:25]
  wire [3:0] _GEN_167 = audioPipeline_io_out_valid ? 4'h7 : stateReg; // @[ChannelController.scala 185:{40,51} 88:25]
  wire [3:0] _stateReg_T_1 = channelCounterWrap ? 4'h9 : 4'h2; // @[ChannelController.scala 192:37]
  wire [3:0] _GEN_168 = outputCounterWrap_wrap_wrap ? 4'h1 : stateReg; // @[ChannelController.scala 196:{31,42} 88:25]
  wire [3:0] _GEN_169 = 4'h9 == stateReg ? _GEN_168 : stateReg; // @[ChannelController.scala 158:20 88:25]
  wire [3:0] _GEN_170 = 4'h8 == stateReg ? _stateReg_T_1 : _GEN_169; // @[ChannelController.scala 158:20 192:31]
  wire [3:0] _GEN_171 = 4'h7 == stateReg ? 4'h8 : _GEN_170; // @[ChannelController.scala 158:20 189:32]
  wire [3:0] _GEN_172 = 4'h6 == stateReg ? _GEN_167 : _GEN_171; // @[ChannelController.scala 158:20]
  wire [3:0] _GEN_173 = 4'h5 == stateReg ? _GEN_166 : _GEN_172; // @[ChannelController.scala 158:20]
  wire [3:0] _GEN_174 = 4'h4 == stateReg ? _stateReg_T : _GEN_173; // @[ChannelController.scala 158:20 176:32]
  wire [3:0] _GEN_175 = 4'h3 == stateReg ? 4'h4 : _GEN_174; // @[ChannelController.scala 158:20 173:32]
  wire [16:0] _io_audio_bits_T_1 = $signed(accumulatorReg_left) < -17'sh8000 ? $signed(-17'sh8000) : $signed(
    accumulatorReg_left); // @[Util.scala 264:51]
  wire [16:0] io_audio_bits_sample_left = $signed(_io_audio_bits_T_1) < 17'sh7fff ? $signed(_io_audio_bits_T_1) :
    $signed(17'sh7fff); // @[Util.scala 264:60]
  AudioPipeline audioPipeline ( // @[ChannelController.scala 104:29]
    .clock(audioPipeline_clock),
    .reset(audioPipeline_reset),
    .io_in_ready(audioPipeline_io_in_ready),
    .io_in_valid(audioPipeline_io_in_valid),
    .io_in_bits_state_samples_0(audioPipeline_io_in_bits_state_samples_0),
    .io_in_bits_state_samples_1(audioPipeline_io_in_bits_state_samples_1),
    .io_in_bits_state_underflow(audioPipeline_io_in_bits_state_underflow),
    .io_in_bits_state_adpcmStep(audioPipeline_io_in_bits_state_adpcmStep),
    .io_in_bits_state_lerpIndex(audioPipeline_io_in_bits_state_lerpIndex),
    .io_in_bits_state_loopEnable(audioPipeline_io_in_bits_state_loopEnable),
    .io_in_bits_state_loopStep(audioPipeline_io_in_bits_state_loopStep),
    .io_in_bits_state_loopSample(audioPipeline_io_in_bits_state_loopSample),
    .io_in_bits_pitch(audioPipeline_io_in_bits_pitch),
    .io_in_bits_level(audioPipeline_io_in_bits_level),
    .io_in_bits_pan(audioPipeline_io_in_bits_pan),
    .io_out_valid(audioPipeline_io_out_valid),
    .io_out_bits_state_samples_0(audioPipeline_io_out_bits_state_samples_0),
    .io_out_bits_state_samples_1(audioPipeline_io_out_bits_state_samples_1),
    .io_out_bits_state_underflow(audioPipeline_io_out_bits_state_underflow),
    .io_out_bits_state_adpcmStep(audioPipeline_io_out_bits_state_adpcmStep),
    .io_out_bits_state_lerpIndex(audioPipeline_io_out_bits_state_lerpIndex),
    .io_out_bits_state_loopEnable(audioPipeline_io_out_bits_state_loopEnable),
    .io_out_bits_state_loopStep(audioPipeline_io_out_bits_state_loopStep),
    .io_out_bits_state_loopSample(audioPipeline_io_out_bits_state_loopSample),
    .io_out_bits_audio_left(audioPipeline_io_out_bits_audio_left),
    .io_pcmData_ready(audioPipeline_io_pcmData_ready),
    .io_pcmData_valid(audioPipeline_io_pcmData_valid),
    .io_pcmData_bits(audioPipeline_io_pcmData_bits),
    .io_loopStart(audioPipeline_io_loopStart)
  );
  assign channelStateMem_channelState_MPORT_en = channelStateMem_channelState_MPORT_en_pipe_0;
  assign channelStateMem_channelState_MPORT_addr = channelStateMem_channelState_MPORT_addr_pipe_0;
  assign channelStateMem_channelState_MPORT_data = channelStateMem[channelStateMem_channelState_MPORT_addr]; // @[ChannelController.scala 99:36]
  assign channelStateMem_MPORT_data = {hi,lo};
  assign channelStateMem_MPORT_addr = channelCounter;
  assign channelStateMem_MPORT_mask = 1'h1;
  assign channelStateMem_MPORT_en = _T | _T_10;
  assign io_done = _T_4 & channelStateReg_done; // @[ChannelController.scala 203:39]
  assign io_index = channelCounter; // @[ChannelController.scala 201:12]
  assign io_audio_valid = outputCounterWrap_value == 9'h16a; // @[Counter.scala 45:24]
  assign io_audio_bits_left = io_audio_bits_sample_left[15:0]; // @[ChannelController.scala 205:17]
  assign io_rom_rd = audioPipeline_io_pcmData_ready & ~pendingReg; // @[ChannelController.scala 122:48]
  assign io_rom_addr = channelStateReg_addr; // @[ChannelController.scala 207:15]
  assign audioPipeline_clock = clock;
  assign audioPipeline_reset = reset;
  assign audioPipeline_io_in_valid = stateReg == 4'h5; // @[ChannelController.scala 105:41]
  assign audioPipeline_io_in_bits_state_samples_0 = channelStateReg_audioPipelineState_samples_0; // @[ChannelController.scala 106:34]
  assign audioPipeline_io_in_bits_state_samples_1 = channelStateReg_audioPipelineState_samples_1; // @[ChannelController.scala 106:34]
  assign audioPipeline_io_in_bits_state_underflow = channelStateReg_audioPipelineState_underflow; // @[ChannelController.scala 106:34]
  assign audioPipeline_io_in_bits_state_adpcmStep = channelStateReg_audioPipelineState_adpcmStep; // @[ChannelController.scala 106:34]
  assign audioPipeline_io_in_bits_state_lerpIndex = channelStateReg_audioPipelineState_lerpIndex; // @[ChannelController.scala 106:34]
  assign audioPipeline_io_in_bits_state_loopEnable = channelStateReg_audioPipelineState_loopEnable; // @[ChannelController.scala 106:34]
  assign audioPipeline_io_in_bits_state_loopStep = channelStateReg_audioPipelineState_loopStep; // @[ChannelController.scala 106:34]
  assign audioPipeline_io_in_bits_state_loopSample = channelStateReg_audioPipelineState_loopSample; // @[ChannelController.scala 106:34]
  assign audioPipeline_io_in_bits_pitch = 3'h7 == channelCounter ? io_regs_7_pitch : _GEN_33; // @[ChannelController.scala 107:{34,34}]
  assign audioPipeline_io_in_bits_level = 3'h7 == channelCounter ? io_regs_7_level : _GEN_41; // @[ChannelController.scala 108:{34,34}]
  assign audioPipeline_io_in_bits_pan = 3'h7 == channelCounter ? io_regs_7_pan : _GEN_49; // @[ChannelController.scala 109:{32,32}]
  assign audioPipeline_io_pcmData_valid = io_rom_valid; // @[ChannelController.scala 110:34]
  assign audioPipeline_io_pcmData_bits = channelStateReg_nibble ? io_rom_dout[3:0] : io_rom_dout[7:4]; // @[ChannelController.scala 111:39]
  assign audioPipeline_io_loopStart = channelStateReg_loopStart; // @[ChannelController.scala 112:30]
  always @(posedge clock) begin
    if (channelStateMem_MPORT_en & channelStateMem_MPORT_mask) begin
      channelStateMem[channelStateMem_MPORT_addr] <= channelStateMem_MPORT_data; // @[ChannelController.scala 99:36]
    end
    channelStateMem_channelState_MPORT_en_pipe_0 <= stateReg == 4'h2;
    if (stateReg == 4'h2) begin
      channelStateMem_channelState_MPORT_addr_pipe_0 <= channelCounter;
    end
    if (reset) begin // @[ChannelController.scala 88:25]
      stateReg <= 4'h0; // @[ChannelController.scala 88:25]
    end else if (4'h0 == stateReg) begin // @[ChannelController.scala 158:20]
      if (channelCounterWrap) begin // @[ChannelController.scala 161:32]
        stateReg <= 4'h1; // @[ChannelController.scala 161:43]
      end
    end else if (4'h1 == stateReg) begin // @[ChannelController.scala 158:20]
      if (io_enable) begin // @[ChannelController.scala 166:23]
        stateReg <= 4'h2; // @[ChannelController.scala 166:34]
      end
    end else if (4'h2 == stateReg) begin // @[ChannelController.scala 158:20]
      stateReg <= 4'h3; // @[ChannelController.scala 170:31]
    end else begin
      stateReg <= _GEN_175;
    end
    if (audioPipeline_io_out_valid) begin // @[ChannelController.scala 143:36]
      accumulatorReg_left <= accumulatorReg_sample_1_left; // @[ChannelController.scala 145:20]
    end else if (stateReg == 4'h1) begin // @[ChannelController.scala 126:33]
      accumulatorReg_left <= 17'sh0; // @[ChannelController.scala 126:50]
    end
    if (reset) begin // @[Counter.scala 40:34]
      channelCounter <= 3'h0; // @[Counter.scala 40:34]
    end else if (_T_2) begin // @[Counter.scala 86:48]
      channelCounter <= _wrap_value_T_1; // @[Counter.scala 46:13]
    end
    if (reset) begin // @[Counter.scala 40:34]
      outputCounterWrap_value <= 9'h0; // @[Counter.scala 40:34]
    end else if (outputCounterWrap_wrap_wrap) begin // @[Counter.scala 48:20]
      outputCounterWrap_value <= 9'h0; // @[Counter.scala 48:28]
    end else begin
      outputCounterWrap_value <= _outputCounterWrap_wrap_value_T_1; // @[Counter.scala 46:13]
    end
    if (stateReg == 4'h4) begin // @[ChannelController.scala 129:34]
      channelStateReg_enable <= _GEN_75;
    end else if (_channelStateReg_T) begin // @[Reg.scala 20:18]
      channelStateReg_enable <= channelState_enable; // @[Reg.scala 20:22]
    end
    if (_T_5) begin // @[ChannelController.scala 140:39]
      if (channelStateReg_nibble) begin // @[ChannelState.scala 83:18]
        if (_GEN_118 & channelStateReg_addr == _GEN_126) begin // @[ChannelState.scala 84:70]
          channelStateReg_active <= _GEN_90;
        end else if (channelStateReg_addr == _GEN_134) begin // @[ChannelState.scala 86:47]
          channelStateReg_active <= 1'h0; // @[ChannelState.scala 87:16]
        end else begin
          channelStateReg_active <= _GEN_90;
        end
      end else begin
        channelStateReg_active <= _GEN_90;
      end
    end else begin
      channelStateReg_active <= _GEN_90;
    end
    if (_T_5) begin // @[ChannelController.scala 140:39]
      if (channelStateReg_nibble) begin // @[ChannelState.scala 83:18]
        if (_GEN_118 & channelStateReg_addr == _GEN_126) begin // @[ChannelState.scala 84:70]
          channelStateReg_done <= _GEN_91;
        end else begin
          channelStateReg_done <= _GEN_136;
        end
      end else begin
        channelStateReg_done <= _GEN_91;
      end
    end else begin
      channelStateReg_done <= _GEN_91;
    end
    if (_T_5) begin // @[ChannelController.scala 140:39]
      channelStateReg_nibble <= _channelStateReg_loopStart_T_2; // @[ChannelState.scala 82:12]
    end else if (stateReg == 4'h4) begin // @[ChannelController.scala 129:34]
      if (start) begin // @[ChannelController.scala 130:17]
        channelStateReg_nibble <= 1'h0; // @[ChannelState.scala 60:12]
      end else begin
        channelStateReg_nibble <= _GEN_16;
      end
    end else begin
      channelStateReg_nibble <= _GEN_16;
    end
    if (_T_5) begin // @[ChannelController.scala 140:39]
      if (channelStateReg_nibble) begin // @[ChannelState.scala 83:18]
        if (_GEN_118 & channelStateReg_addr == _GEN_126) begin // @[ChannelState.scala 84:70]
          if (3'h7 == channelCounter) begin // @[ChannelState.scala 81:48]
            channelStateReg_addr <= io_regs_7_loopStartAddr; // @[ChannelState.scala 81:48]
          end else begin
            channelStateReg_addr <= _GEN_109;
          end
        end else if (channelStateReg_addr == _GEN_134) begin // @[ChannelState.scala 86:47]
          channelStateReg_addr <= _GEN_93;
        end else begin
          channelStateReg_addr <= _channelStateReg_addr_T_1; // @[ChannelState.scala 90:14]
        end
      end else begin
        channelStateReg_addr <= _GEN_93;
      end
    end else begin
      channelStateReg_addr <= _GEN_93;
    end
    if (_T_5) begin // @[ChannelController.scala 140:39]
      channelStateReg_loopStart <= _GEN_118 & channelStateReg_addr == _GEN_110 & ~channelStateReg_nibble; // @[ChannelState.scala 81:15]
    end else if (stateReg == 4'h4) begin // @[ChannelController.scala 129:34]
      if (start) begin // @[ChannelController.scala 130:17]
        channelStateReg_loopStart <= 1'h0; // @[ChannelState.scala 62:15]
      end else begin
        channelStateReg_loopStart <= _GEN_18;
      end
    end else begin
      channelStateReg_loopStart <= _GEN_18;
    end
    if (audioPipeline_io_out_valid) begin // @[ChannelController.scala 143:36]
      channelStateReg_audioPipelineState_samples_0 <= audioPipeline_io_out_bits_state_samples_0; // @[ChannelController.scala 148:40]
    end else if (stateReg == 4'h4) begin // @[ChannelController.scala 129:34]
      if (start) begin // @[ChannelController.scala 130:17]
        channelStateReg_audioPipelineState_samples_0 <= 16'sh0; // @[ChannelState.scala 63:24]
      end else begin
        channelStateReg_audioPipelineState_samples_0 <= _GEN_19;
      end
    end else begin
      channelStateReg_audioPipelineState_samples_0 <= _GEN_19;
    end
    if (audioPipeline_io_out_valid) begin // @[ChannelController.scala 143:36]
      channelStateReg_audioPipelineState_samples_1 <= audioPipeline_io_out_bits_state_samples_1; // @[ChannelController.scala 148:40]
    end else if (stateReg == 4'h4) begin // @[ChannelController.scala 129:34]
      if (start) begin // @[ChannelController.scala 130:17]
        channelStateReg_audioPipelineState_samples_1 <= 16'sh0; // @[ChannelState.scala 63:24]
      end else begin
        channelStateReg_audioPipelineState_samples_1 <= _GEN_20;
      end
    end else begin
      channelStateReg_audioPipelineState_samples_1 <= _GEN_20;
    end
    if (audioPipeline_io_out_valid) begin // @[ChannelController.scala 143:36]
      channelStateReg_audioPipelineState_underflow <= audioPipeline_io_out_bits_state_underflow; // @[ChannelController.scala 148:40]
    end else if (stateReg == 4'h4) begin // @[ChannelController.scala 129:34]
      channelStateReg_audioPipelineState_underflow <= _GEN_83;
    end else if (_channelStateReg_T) begin // @[Reg.scala 20:18]
      channelStateReg_audioPipelineState_underflow <= channelState_audioPipelineState_underflow; // @[Reg.scala 20:22]
    end
    if (audioPipeline_io_out_valid) begin // @[ChannelController.scala 143:36]
      channelStateReg_audioPipelineState_adpcmStep <= audioPipeline_io_out_bits_state_adpcmStep; // @[ChannelController.scala 148:40]
    end else if (stateReg == 4'h4) begin // @[ChannelController.scala 129:34]
      if (start) begin // @[ChannelController.scala 130:17]
        channelStateReg_audioPipelineState_adpcmStep <= 16'sh7f; // @[ChannelState.scala 63:24]
      end else begin
        channelStateReg_audioPipelineState_adpcmStep <= _GEN_22;
      end
    end else begin
      channelStateReg_audioPipelineState_adpcmStep <= _GEN_22;
    end
    if (audioPipeline_io_out_valid) begin // @[ChannelController.scala 143:36]
      channelStateReg_audioPipelineState_lerpIndex <= audioPipeline_io_out_bits_state_lerpIndex; // @[ChannelController.scala 148:40]
    end else if (stateReg == 4'h4) begin // @[ChannelController.scala 129:34]
      if (start) begin // @[ChannelController.scala 130:17]
        channelStateReg_audioPipelineState_lerpIndex <= 10'h0; // @[ChannelState.scala 63:24]
      end else begin
        channelStateReg_audioPipelineState_lerpIndex <= _GEN_23;
      end
    end else begin
      channelStateReg_audioPipelineState_lerpIndex <= _GEN_23;
    end
    if (audioPipeline_io_out_valid) begin // @[ChannelController.scala 143:36]
      channelStateReg_audioPipelineState_loopEnable <= audioPipeline_io_out_bits_state_loopEnable; // @[ChannelController.scala 148:40]
    end else if (stateReg == 4'h4) begin // @[ChannelController.scala 129:34]
      if (start) begin // @[ChannelController.scala 130:17]
        channelStateReg_audioPipelineState_loopEnable <= 1'h0; // @[ChannelState.scala 63:24]
      end else begin
        channelStateReg_audioPipelineState_loopEnable <= _GEN_24;
      end
    end else begin
      channelStateReg_audioPipelineState_loopEnable <= _GEN_24;
    end
    if (audioPipeline_io_out_valid) begin // @[ChannelController.scala 143:36]
      channelStateReg_audioPipelineState_loopStep <= audioPipeline_io_out_bits_state_loopStep; // @[ChannelController.scala 148:40]
    end else if (stateReg == 4'h4) begin // @[ChannelController.scala 129:34]
      if (start) begin // @[ChannelController.scala 130:17]
        channelStateReg_audioPipelineState_loopStep <= 16'sh0; // @[ChannelState.scala 63:24]
      end else begin
        channelStateReg_audioPipelineState_loopStep <= _GEN_25;
      end
    end else begin
      channelStateReg_audioPipelineState_loopStep <= _GEN_25;
    end
    if (audioPipeline_io_out_valid) begin // @[ChannelController.scala 143:36]
      channelStateReg_audioPipelineState_loopSample <= audioPipeline_io_out_bits_state_loopSample; // @[ChannelController.scala 148:40]
    end else if (stateReg == 4'h4) begin // @[ChannelController.scala 129:34]
      if (start) begin // @[ChannelController.scala 130:17]
        channelStateReg_audioPipelineState_loopSample <= 16'sh0; // @[ChannelState.scala 63:24]
      end else begin
        channelStateReg_audioPipelineState_loopSample <= _GEN_26;
      end
    end else begin
      channelStateReg_audioPipelineState_loopSample <= _GEN_26;
    end
    if (reset) begin // @[Util.scala 218:28]
      pendingReg <= 1'h0; // @[Util.scala 218:28]
    end else if (io_rom_valid) begin // @[Util.scala 219:17]
      pendingReg <= 1'h0; // @[Util.scala 219:29]
    end else begin
      pendingReg <= _GEN_59;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    channelStateMem[initvar] = _RAND_0[120:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  channelStateMem_channelState_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  channelStateMem_channelState_MPORT_addr_pipe_0 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  stateReg = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  accumulatorReg_left = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  channelCounter = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  outputCounterWrap_value = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  channelStateReg_enable = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  channelStateReg_active = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  channelStateReg_done = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  channelStateReg_nibble = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  channelStateReg_addr = _RAND_11[23:0];
  _RAND_12 = {1{`RANDOM}};
  channelStateReg_loopStart = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  channelStateReg_audioPipelineState_samples_0 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  channelStateReg_audioPipelineState_samples_1 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  channelStateReg_audioPipelineState_underflow = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  channelStateReg_audioPipelineState_adpcmStep = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  channelStateReg_audioPipelineState_lerpIndex = _RAND_17[9:0];
  _RAND_18 = {1{`RANDOM}};
  channelStateReg_audioPipelineState_loopEnable = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  channelStateReg_audioPipelineState_loopStep = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  channelStateReg_audioPipelineState_loopSample = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  pendingReg = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module YMZ280B(
  input         clock,
  input         reset,
  input         io_cpu_rd,
  input         io_cpu_wr,
  input         io_cpu_addr,
  input  [7:0]  io_cpu_din,
  output [7:0]  io_cpu_dout,
  output        io_rom_rd,
  output [23:0] io_rom_addr,
  input  [7:0]  io_rom_dout,
  input         io_rom_wait_n,
  input         io_rom_valid,
  output        io_audio_valid,
  output [15:0] io_audio_bits_left,
  output        io_irq
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
`endif // RANDOMIZE_REG_INIT
  wire  channelCtrl_clock; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_reset; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_0_pitch; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_0_flags_keyOn; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_0_flags_loop; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_0_level; // @[YMZ280B.scala 117:27]
  wire [3:0] channelCtrl_io_regs_0_pan; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_0_startAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_0_loopStartAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_0_loopEndAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_0_endAddr; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_1_pitch; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_1_flags_keyOn; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_1_flags_loop; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_1_level; // @[YMZ280B.scala 117:27]
  wire [3:0] channelCtrl_io_regs_1_pan; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_1_startAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_1_loopStartAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_1_loopEndAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_1_endAddr; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_2_pitch; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_2_flags_keyOn; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_2_flags_loop; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_2_level; // @[YMZ280B.scala 117:27]
  wire [3:0] channelCtrl_io_regs_2_pan; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_2_startAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_2_loopStartAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_2_loopEndAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_2_endAddr; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_3_pitch; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_3_flags_keyOn; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_3_flags_loop; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_3_level; // @[YMZ280B.scala 117:27]
  wire [3:0] channelCtrl_io_regs_3_pan; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_3_startAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_3_loopStartAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_3_loopEndAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_3_endAddr; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_4_pitch; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_4_flags_keyOn; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_4_flags_loop; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_4_level; // @[YMZ280B.scala 117:27]
  wire [3:0] channelCtrl_io_regs_4_pan; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_4_startAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_4_loopStartAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_4_loopEndAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_4_endAddr; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_5_pitch; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_5_flags_keyOn; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_5_flags_loop; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_5_level; // @[YMZ280B.scala 117:27]
  wire [3:0] channelCtrl_io_regs_5_pan; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_5_startAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_5_loopStartAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_5_loopEndAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_5_endAddr; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_6_pitch; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_6_flags_keyOn; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_6_flags_loop; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_6_level; // @[YMZ280B.scala 117:27]
  wire [3:0] channelCtrl_io_regs_6_pan; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_6_startAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_6_loopStartAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_6_loopEndAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_6_endAddr; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_7_pitch; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_7_flags_keyOn; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_regs_7_flags_loop; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_regs_7_level; // @[YMZ280B.scala 117:27]
  wire [3:0] channelCtrl_io_regs_7_pan; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_7_startAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_7_loopStartAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_7_loopEndAddr; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_regs_7_endAddr; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_enable; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_done; // @[YMZ280B.scala 117:27]
  wire [2:0] channelCtrl_io_index; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_audio_valid; // @[YMZ280B.scala 117:27]
  wire [15:0] channelCtrl_io_audio_bits_left; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_rom_rd; // @[YMZ280B.scala 117:27]
  wire [23:0] channelCtrl_io_rom_addr; // @[YMZ280B.scala 117:27]
  wire [7:0] channelCtrl_io_rom_dout; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_rom_wait_n; // @[YMZ280B.scala 117:27]
  wire  channelCtrl_io_rom_valid; // @[YMZ280B.scala 117:27]
  reg [7:0] addrReg; // @[YMZ280B.scala 105:24]
  reg [7:0] dataReg; // @[YMZ280B.scala 106:24]
  reg [7:0] statusReg; // @[YMZ280B.scala 107:26]
  reg [7:0] registerFile_0; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_1; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_2; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_3; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_4; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_5; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_6; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_7; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_8; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_9; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_10; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_11; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_12; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_13; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_14; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_15; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_16; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_17; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_18; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_19; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_20; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_21; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_22; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_23; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_24; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_25; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_26; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_27; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_28; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_29; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_30; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_31; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_32; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_33; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_34; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_35; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_36; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_37; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_38; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_39; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_40; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_41; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_42; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_43; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_44; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_45; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_46; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_47; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_48; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_49; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_50; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_51; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_52; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_53; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_54; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_55; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_56; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_57; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_58; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_59; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_60; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_61; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_62; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_63; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_64; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_65; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_66; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_67; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_68; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_69; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_70; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_71; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_72; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_73; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_74; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_75; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_76; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_77; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_78; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_79; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_80; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_81; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_82; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_83; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_84; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_85; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_86; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_87; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_88; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_89; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_90; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_91; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_92; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_93; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_94; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_95; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_96; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_97; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_98; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_99; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_100; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_101; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_102; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_103; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_104; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_105; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_106; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_107; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_108; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_109; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_110; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_111; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_112; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_113; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_114; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_115; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_116; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_117; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_118; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_119; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_120; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_121; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_122; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_123; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_124; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_125; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_126; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_127; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_254; // @[YMZ280B.scala 108:29]
  reg [7:0] registerFile_255; // @[YMZ280B.scala 108:29]
  wire [63:0] channelRegs_lo = {registerFile_65,registerFile_97,registerFile_34,registerFile_66,registerFile_98,
    registerFile_35,registerFile_67,registerFile_99}; // @[Cat.scala 33:92]
  wire [119:0] _channelRegs_T_2 = {registerFile_0,registerFile_1[7:4],registerFile_2,registerFile_3[3:0],registerFile_32
    ,registerFile_64,registerFile_96,registerFile_33,channelRegs_lo}; // @[Cat.scala 33:92]
  wire [63:0] channelRegs_lo_1 = {registerFile_69,registerFile_101,registerFile_38,registerFile_70,registerFile_102,
    registerFile_39,registerFile_71,registerFile_103}; // @[Cat.scala 33:92]
  wire [119:0] _channelRegs_T_15 = {registerFile_4,registerFile_5[7:4],registerFile_6,registerFile_7[3:0],
    registerFile_36,registerFile_68,registerFile_100,registerFile_37,channelRegs_lo_1}; // @[Cat.scala 33:92]
  wire [63:0] channelRegs_lo_2 = {registerFile_73,registerFile_105,registerFile_42,registerFile_74,registerFile_106,
    registerFile_43,registerFile_75,registerFile_107}; // @[Cat.scala 33:92]
  wire [119:0] _channelRegs_T_28 = {registerFile_8,registerFile_9[7:4],registerFile_10,registerFile_11[3:0],
    registerFile_40,registerFile_72,registerFile_104,registerFile_41,channelRegs_lo_2}; // @[Cat.scala 33:92]
  wire [63:0] channelRegs_lo_3 = {registerFile_77,registerFile_109,registerFile_46,registerFile_78,registerFile_110,
    registerFile_47,registerFile_79,registerFile_111}; // @[Cat.scala 33:92]
  wire [119:0] _channelRegs_T_41 = {registerFile_12,registerFile_13[7:4],registerFile_14,registerFile_15[3:0],
    registerFile_44,registerFile_76,registerFile_108,registerFile_45,channelRegs_lo_3}; // @[Cat.scala 33:92]
  wire [63:0] channelRegs_lo_4 = {registerFile_81,registerFile_113,registerFile_50,registerFile_82,registerFile_114,
    registerFile_51,registerFile_83,registerFile_115}; // @[Cat.scala 33:92]
  wire [119:0] _channelRegs_T_54 = {registerFile_16,registerFile_17[7:4],registerFile_18,registerFile_19[3:0],
    registerFile_48,registerFile_80,registerFile_112,registerFile_49,channelRegs_lo_4}; // @[Cat.scala 33:92]
  wire [63:0] channelRegs_lo_5 = {registerFile_85,registerFile_117,registerFile_54,registerFile_86,registerFile_118,
    registerFile_55,registerFile_87,registerFile_119}; // @[Cat.scala 33:92]
  wire [119:0] _channelRegs_T_67 = {registerFile_20,registerFile_21[7:4],registerFile_22,registerFile_23[3:0],
    registerFile_52,registerFile_84,registerFile_116,registerFile_53,channelRegs_lo_5}; // @[Cat.scala 33:92]
  wire [63:0] channelRegs_lo_6 = {registerFile_89,registerFile_121,registerFile_58,registerFile_90,registerFile_122,
    registerFile_59,registerFile_91,registerFile_123}; // @[Cat.scala 33:92]
  wire [119:0] _channelRegs_T_80 = {registerFile_24,registerFile_25[7:4],registerFile_26,registerFile_27[3:0],
    registerFile_56,registerFile_88,registerFile_120,registerFile_57,channelRegs_lo_6}; // @[Cat.scala 33:92]
  wire [63:0] channelRegs_lo_7 = {registerFile_93,registerFile_125,registerFile_62,registerFile_94,registerFile_126,
    registerFile_63,registerFile_95,registerFile_127}; // @[Cat.scala 33:92]
  wire [119:0] _channelRegs_T_93 = {registerFile_28,registerFile_29[7:4],registerFile_30,registerFile_31[3:0],
    registerFile_60,registerFile_92,registerFile_124,registerFile_61,channelRegs_lo_7}; // @[Cat.scala 33:92]
  wire [10:0] _utilReg_T_3 = {registerFile_254,registerFile_255[7],registerFile_255[6],registerFile_255[4]}; // @[Cat.scala 33:92]
  wire  utilReg_flags_irqEnable = _utilReg_T_3[0]; // @[UtilReg.scala 65:15]
  wire [7:0] utilReg_irqMask = _utilReg_T_3[10:3]; // @[UtilReg.scala 65:15]
  wire  writeAddr = io_cpu_wr & ~io_cpu_addr; // @[YMZ280B.scala 124:29]
  wire  writeData = io_cpu_wr & io_cpu_addr; // @[YMZ280B.scala 125:29]
  wire  readStatus = io_cpu_rd & io_cpu_addr; // @[YMZ280B.scala 126:30]
  wire [7:0] _statusReg_T = 8'h1 << channelCtrl_io_index; // @[YMZ280B.scala 135:60]
  wire [7:0] _statusReg_T_1 = statusReg | _statusReg_T; // @[YMZ280B.scala 135:60]
  wire [7:0] _io_irq_T = statusReg & utilReg_irqMask; // @[YMZ280B.scala 145:51]
  ChannelController channelCtrl ( // @[YMZ280B.scala 117:27]
    .clock(channelCtrl_clock),
    .reset(channelCtrl_reset),
    .io_regs_0_pitch(channelCtrl_io_regs_0_pitch),
    .io_regs_0_flags_keyOn(channelCtrl_io_regs_0_flags_keyOn),
    .io_regs_0_flags_loop(channelCtrl_io_regs_0_flags_loop),
    .io_regs_0_level(channelCtrl_io_regs_0_level),
    .io_regs_0_pan(channelCtrl_io_regs_0_pan),
    .io_regs_0_startAddr(channelCtrl_io_regs_0_startAddr),
    .io_regs_0_loopStartAddr(channelCtrl_io_regs_0_loopStartAddr),
    .io_regs_0_loopEndAddr(channelCtrl_io_regs_0_loopEndAddr),
    .io_regs_0_endAddr(channelCtrl_io_regs_0_endAddr),
    .io_regs_1_pitch(channelCtrl_io_regs_1_pitch),
    .io_regs_1_flags_keyOn(channelCtrl_io_regs_1_flags_keyOn),
    .io_regs_1_flags_loop(channelCtrl_io_regs_1_flags_loop),
    .io_regs_1_level(channelCtrl_io_regs_1_level),
    .io_regs_1_pan(channelCtrl_io_regs_1_pan),
    .io_regs_1_startAddr(channelCtrl_io_regs_1_startAddr),
    .io_regs_1_loopStartAddr(channelCtrl_io_regs_1_loopStartAddr),
    .io_regs_1_loopEndAddr(channelCtrl_io_regs_1_loopEndAddr),
    .io_regs_1_endAddr(channelCtrl_io_regs_1_endAddr),
    .io_regs_2_pitch(channelCtrl_io_regs_2_pitch),
    .io_regs_2_flags_keyOn(channelCtrl_io_regs_2_flags_keyOn),
    .io_regs_2_flags_loop(channelCtrl_io_regs_2_flags_loop),
    .io_regs_2_level(channelCtrl_io_regs_2_level),
    .io_regs_2_pan(channelCtrl_io_regs_2_pan),
    .io_regs_2_startAddr(channelCtrl_io_regs_2_startAddr),
    .io_regs_2_loopStartAddr(channelCtrl_io_regs_2_loopStartAddr),
    .io_regs_2_loopEndAddr(channelCtrl_io_regs_2_loopEndAddr),
    .io_regs_2_endAddr(channelCtrl_io_regs_2_endAddr),
    .io_regs_3_pitch(channelCtrl_io_regs_3_pitch),
    .io_regs_3_flags_keyOn(channelCtrl_io_regs_3_flags_keyOn),
    .io_regs_3_flags_loop(channelCtrl_io_regs_3_flags_loop),
    .io_regs_3_level(channelCtrl_io_regs_3_level),
    .io_regs_3_pan(channelCtrl_io_regs_3_pan),
    .io_regs_3_startAddr(channelCtrl_io_regs_3_startAddr),
    .io_regs_3_loopStartAddr(channelCtrl_io_regs_3_loopStartAddr),
    .io_regs_3_loopEndAddr(channelCtrl_io_regs_3_loopEndAddr),
    .io_regs_3_endAddr(channelCtrl_io_regs_3_endAddr),
    .io_regs_4_pitch(channelCtrl_io_regs_4_pitch),
    .io_regs_4_flags_keyOn(channelCtrl_io_regs_4_flags_keyOn),
    .io_regs_4_flags_loop(channelCtrl_io_regs_4_flags_loop),
    .io_regs_4_level(channelCtrl_io_regs_4_level),
    .io_regs_4_pan(channelCtrl_io_regs_4_pan),
    .io_regs_4_startAddr(channelCtrl_io_regs_4_startAddr),
    .io_regs_4_loopStartAddr(channelCtrl_io_regs_4_loopStartAddr),
    .io_regs_4_loopEndAddr(channelCtrl_io_regs_4_loopEndAddr),
    .io_regs_4_endAddr(channelCtrl_io_regs_4_endAddr),
    .io_regs_5_pitch(channelCtrl_io_regs_5_pitch),
    .io_regs_5_flags_keyOn(channelCtrl_io_regs_5_flags_keyOn),
    .io_regs_5_flags_loop(channelCtrl_io_regs_5_flags_loop),
    .io_regs_5_level(channelCtrl_io_regs_5_level),
    .io_regs_5_pan(channelCtrl_io_regs_5_pan),
    .io_regs_5_startAddr(channelCtrl_io_regs_5_startAddr),
    .io_regs_5_loopStartAddr(channelCtrl_io_regs_5_loopStartAddr),
    .io_regs_5_loopEndAddr(channelCtrl_io_regs_5_loopEndAddr),
    .io_regs_5_endAddr(channelCtrl_io_regs_5_endAddr),
    .io_regs_6_pitch(channelCtrl_io_regs_6_pitch),
    .io_regs_6_flags_keyOn(channelCtrl_io_regs_6_flags_keyOn),
    .io_regs_6_flags_loop(channelCtrl_io_regs_6_flags_loop),
    .io_regs_6_level(channelCtrl_io_regs_6_level),
    .io_regs_6_pan(channelCtrl_io_regs_6_pan),
    .io_regs_6_startAddr(channelCtrl_io_regs_6_startAddr),
    .io_regs_6_loopStartAddr(channelCtrl_io_regs_6_loopStartAddr),
    .io_regs_6_loopEndAddr(channelCtrl_io_regs_6_loopEndAddr),
    .io_regs_6_endAddr(channelCtrl_io_regs_6_endAddr),
    .io_regs_7_pitch(channelCtrl_io_regs_7_pitch),
    .io_regs_7_flags_keyOn(channelCtrl_io_regs_7_flags_keyOn),
    .io_regs_7_flags_loop(channelCtrl_io_regs_7_flags_loop),
    .io_regs_7_level(channelCtrl_io_regs_7_level),
    .io_regs_7_pan(channelCtrl_io_regs_7_pan),
    .io_regs_7_startAddr(channelCtrl_io_regs_7_startAddr),
    .io_regs_7_loopStartAddr(channelCtrl_io_regs_7_loopStartAddr),
    .io_regs_7_loopEndAddr(channelCtrl_io_regs_7_loopEndAddr),
    .io_regs_7_endAddr(channelCtrl_io_regs_7_endAddr),
    .io_enable(channelCtrl_io_enable),
    .io_done(channelCtrl_io_done),
    .io_index(channelCtrl_io_index),
    .io_audio_valid(channelCtrl_io_audio_valid),
    .io_audio_bits_left(channelCtrl_io_audio_bits_left),
    .io_rom_rd(channelCtrl_io_rom_rd),
    .io_rom_addr(channelCtrl_io_rom_addr),
    .io_rom_dout(channelCtrl_io_rom_dout),
    .io_rom_wait_n(channelCtrl_io_rom_wait_n),
    .io_rom_valid(channelCtrl_io_rom_valid)
  );
  assign io_cpu_dout = dataReg; // @[YMZ280B.scala 144:15]
  assign io_rom_rd = channelCtrl_io_rom_rd; // @[YMZ280B.scala 121:22]
  assign io_rom_addr = channelCtrl_io_rom_addr; // @[YMZ280B.scala 121:22]
  assign io_audio_valid = channelCtrl_io_audio_valid; // @[YMZ280B.scala 120:24]
  assign io_audio_bits_left = channelCtrl_io_audio_bits_left; // @[YMZ280B.scala 120:24]
  assign io_irq = utilReg_flags_irqEnable & |_io_irq_T; // @[YMZ280B.scala 145:37]
  assign channelCtrl_clock = clock;
  assign channelCtrl_reset = reset;
  assign channelCtrl_io_regs_0_pitch = _channelRegs_T_2[119:112]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_0_flags_keyOn = _channelRegs_T_2[111]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_0_flags_loop = _channelRegs_T_2[108]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_0_level = _channelRegs_T_2[107:100]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_0_pan = _channelRegs_T_2[99:96]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_0_startAddr = _channelRegs_T_2[95:72]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_0_loopStartAddr = _channelRegs_T_2[71:48]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_0_loopEndAddr = _channelRegs_T_2[47:24]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_0_endAddr = _channelRegs_T_2[23:0]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_1_pitch = _channelRegs_T_15[119:112]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_1_flags_keyOn = _channelRegs_T_15[111]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_1_flags_loop = _channelRegs_T_15[108]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_1_level = _channelRegs_T_15[107:100]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_1_pan = _channelRegs_T_15[99:96]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_1_startAddr = _channelRegs_T_15[95:72]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_1_loopStartAddr = _channelRegs_T_15[71:48]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_1_loopEndAddr = _channelRegs_T_15[47:24]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_1_endAddr = _channelRegs_T_15[23:0]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_2_pitch = _channelRegs_T_28[119:112]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_2_flags_keyOn = _channelRegs_T_28[111]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_2_flags_loop = _channelRegs_T_28[108]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_2_level = _channelRegs_T_28[107:100]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_2_pan = _channelRegs_T_28[99:96]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_2_startAddr = _channelRegs_T_28[95:72]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_2_loopStartAddr = _channelRegs_T_28[71:48]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_2_loopEndAddr = _channelRegs_T_28[47:24]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_2_endAddr = _channelRegs_T_28[23:0]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_3_pitch = _channelRegs_T_41[119:112]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_3_flags_keyOn = _channelRegs_T_41[111]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_3_flags_loop = _channelRegs_T_41[108]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_3_level = _channelRegs_T_41[107:100]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_3_pan = _channelRegs_T_41[99:96]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_3_startAddr = _channelRegs_T_41[95:72]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_3_loopStartAddr = _channelRegs_T_41[71:48]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_3_loopEndAddr = _channelRegs_T_41[47:24]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_3_endAddr = _channelRegs_T_41[23:0]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_4_pitch = _channelRegs_T_54[119:112]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_4_flags_keyOn = _channelRegs_T_54[111]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_4_flags_loop = _channelRegs_T_54[108]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_4_level = _channelRegs_T_54[107:100]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_4_pan = _channelRegs_T_54[99:96]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_4_startAddr = _channelRegs_T_54[95:72]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_4_loopStartAddr = _channelRegs_T_54[71:48]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_4_loopEndAddr = _channelRegs_T_54[47:24]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_4_endAddr = _channelRegs_T_54[23:0]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_5_pitch = _channelRegs_T_67[119:112]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_5_flags_keyOn = _channelRegs_T_67[111]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_5_flags_loop = _channelRegs_T_67[108]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_5_level = _channelRegs_T_67[107:100]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_5_pan = _channelRegs_T_67[99:96]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_5_startAddr = _channelRegs_T_67[95:72]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_5_loopStartAddr = _channelRegs_T_67[71:48]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_5_loopEndAddr = _channelRegs_T_67[47:24]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_5_endAddr = _channelRegs_T_67[23:0]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_6_pitch = _channelRegs_T_80[119:112]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_6_flags_keyOn = _channelRegs_T_80[111]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_6_flags_loop = _channelRegs_T_80[108]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_6_level = _channelRegs_T_80[107:100]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_6_pan = _channelRegs_T_80[99:96]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_6_startAddr = _channelRegs_T_80[95:72]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_6_loopStartAddr = _channelRegs_T_80[71:48]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_6_loopEndAddr = _channelRegs_T_80[47:24]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_6_endAddr = _channelRegs_T_80[23:0]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_7_pitch = _channelRegs_T_93[119:112]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_7_flags_keyOn = _channelRegs_T_93[111]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_7_flags_loop = _channelRegs_T_93[108]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_7_level = _channelRegs_T_93[107:100]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_7_pan = _channelRegs_T_93[99:96]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_7_startAddr = _channelRegs_T_93[95:72]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_7_loopStartAddr = _channelRegs_T_93[71:48]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_7_loopEndAddr = _channelRegs_T_93[47:24]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_regs_7_endAddr = _channelRegs_T_93[23:0]; // @[ChannelReg.scala 101:15]
  assign channelCtrl_io_enable = _utilReg_T_3[2]; // @[UtilReg.scala 65:15]
  assign channelCtrl_io_rom_dout = io_rom_dout; // @[YMZ280B.scala 121:22]
  assign channelCtrl_io_rom_wait_n = io_rom_wait_n; // @[YMZ280B.scala 121:22]
  assign channelCtrl_io_rom_valid = io_rom_valid; // @[YMZ280B.scala 121:22]
  always @(posedge clock) begin
    if (reset) begin // @[YMZ280B.scala 105:24]
      addrReg <= 8'h0; // @[YMZ280B.scala 105:24]
    end else if (writeAddr) begin // @[YMZ280B.scala 129:19]
      addrReg <= io_cpu_din; // @[YMZ280B.scala 129:29]
    end
    if (reset) begin // @[YMZ280B.scala 106:24]
      dataReg <= 8'h0; // @[YMZ280B.scala 106:24]
    end else if (readStatus) begin // @[YMZ280B.scala 138:20]
      dataReg <= statusReg; // @[YMZ280B.scala 139:13]
    end
    if (reset) begin // @[YMZ280B.scala 107:26]
      statusReg <= 8'h0; // @[YMZ280B.scala 107:26]
    end else if (readStatus) begin // @[YMZ280B.scala 138:20]
      statusReg <= 8'h0; // @[YMZ280B.scala 140:15]
    end else if (channelCtrl_io_done) begin // @[YMZ280B.scala 135:29]
      statusReg <= _statusReg_T_1; // @[YMZ280B.scala 135:41]
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_0 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h0 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_0 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_1 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h1 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_1 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_2 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h2 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_2 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_3 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h3 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_3 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_4 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h4 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_4 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_5 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h5 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_5 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_6 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h6 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_6 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_7 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h7 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_7 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_8 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h8 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_8 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_9 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h9 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_9 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_10 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'ha == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_10 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_11 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'hb == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_11 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_12 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'hc == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_12 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_13 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'hd == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_13 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_14 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'he == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_14 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_15 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'hf == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_15 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_16 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h10 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_16 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_17 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h11 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_17 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_18 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h12 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_18 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_19 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h13 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_19 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_20 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h14 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_20 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_21 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h15 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_21 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_22 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h16 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_22 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_23 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h17 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_23 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_24 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h18 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_24 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_25 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h19 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_25 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_26 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h1a == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_26 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_27 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h1b == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_27 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_28 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h1c == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_28 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_29 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h1d == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_29 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_30 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h1e == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_30 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_31 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h1f == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_31 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_32 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h20 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_32 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_33 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h21 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_33 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_34 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h22 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_34 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_35 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h23 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_35 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_36 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h24 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_36 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_37 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h25 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_37 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_38 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h26 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_38 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_39 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h27 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_39 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_40 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h28 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_40 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_41 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h29 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_41 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_42 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h2a == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_42 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_43 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h2b == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_43 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_44 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h2c == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_44 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_45 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h2d == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_45 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_46 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h2e == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_46 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_47 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h2f == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_47 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_48 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h30 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_48 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_49 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h31 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_49 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_50 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h32 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_50 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_51 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h33 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_51 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_52 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h34 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_52 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_53 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h35 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_53 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_54 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h36 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_54 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_55 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h37 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_55 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_56 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h38 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_56 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_57 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h39 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_57 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_58 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h3a == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_58 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_59 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h3b == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_59 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_60 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h3c == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_60 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_61 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h3d == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_61 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_62 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h3e == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_62 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_63 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h3f == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_63 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_64 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h40 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_64 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_65 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h41 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_65 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_66 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h42 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_66 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_67 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h43 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_67 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_68 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h44 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_68 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_69 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h45 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_69 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_70 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h46 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_70 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_71 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h47 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_71 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_72 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h48 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_72 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_73 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h49 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_73 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_74 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h4a == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_74 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_75 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h4b == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_75 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_76 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h4c == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_76 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_77 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h4d == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_77 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_78 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h4e == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_78 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_79 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h4f == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_79 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_80 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h50 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_80 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_81 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h51 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_81 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_82 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h52 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_82 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_83 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h53 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_83 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_84 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h54 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_84 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_85 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h55 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_85 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_86 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h56 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_86 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_87 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h57 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_87 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_88 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h58 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_88 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_89 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h59 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_89 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_90 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h5a == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_90 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_91 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h5b == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_91 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_92 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h5c == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_92 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_93 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h5d == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_93 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_94 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h5e == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_94 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_95 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h5f == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_95 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_96 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h60 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_96 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_97 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h61 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_97 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_98 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h62 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_98 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_99 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h63 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_99 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_100 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h64 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_100 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_101 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h65 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_101 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_102 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h66 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_102 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_103 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h67 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_103 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_104 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h68 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_104 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_105 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h69 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_105 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_106 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h6a == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_106 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_107 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h6b == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_107 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_108 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h6c == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_108 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_109 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h6d == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_109 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_110 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h6e == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_110 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_111 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h6f == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_111 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_112 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h70 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_112 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_113 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h71 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_113 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_114 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h72 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_114 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_115 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h73 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_115 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_116 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h74 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_116 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_117 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h75 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_117 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_118 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h76 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_118 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_119 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h77 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_119 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_120 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h78 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_120 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_121 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h79 == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_121 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_122 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h7a == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_122 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_123 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h7b == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_123 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_124 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h7c == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_124 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_125 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h7d == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_125 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_126 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h7e == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_126 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_127 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'h7f == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_127 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_254 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'hfe == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_254 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
    if (reset) begin // @[YMZ280B.scala 108:29]
      registerFile_255 <= 8'h0; // @[YMZ280B.scala 108:29]
    end else if (writeData) begin // @[YMZ280B.scala 132:19]
      if (8'hff == addrReg) begin // @[YMZ280B.scala 132:43]
        registerFile_255 <= io_cpu_din; // @[YMZ280B.scala 132:43]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addrReg = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  statusReg = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  registerFile_0 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  registerFile_1 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  registerFile_2 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  registerFile_3 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  registerFile_4 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  registerFile_5 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  registerFile_6 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  registerFile_7 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  registerFile_8 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  registerFile_9 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  registerFile_10 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  registerFile_11 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  registerFile_12 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  registerFile_13 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  registerFile_14 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  registerFile_15 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  registerFile_16 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  registerFile_17 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  registerFile_18 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  registerFile_19 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  registerFile_20 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  registerFile_21 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  registerFile_22 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  registerFile_23 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  registerFile_24 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  registerFile_25 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  registerFile_26 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  registerFile_27 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  registerFile_28 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  registerFile_29 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  registerFile_30 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  registerFile_31 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  registerFile_32 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  registerFile_33 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  registerFile_34 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  registerFile_35 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  registerFile_36 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  registerFile_37 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  registerFile_38 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  registerFile_39 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  registerFile_40 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  registerFile_41 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  registerFile_42 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  registerFile_43 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  registerFile_44 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  registerFile_45 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  registerFile_46 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  registerFile_47 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  registerFile_48 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  registerFile_49 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  registerFile_50 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  registerFile_51 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  registerFile_52 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  registerFile_53 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  registerFile_54 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  registerFile_55 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  registerFile_56 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  registerFile_57 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  registerFile_58 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  registerFile_59 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  registerFile_60 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  registerFile_61 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  registerFile_62 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  registerFile_63 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  registerFile_64 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  registerFile_65 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  registerFile_66 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  registerFile_67 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  registerFile_68 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  registerFile_69 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  registerFile_70 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  registerFile_71 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  registerFile_72 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  registerFile_73 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  registerFile_74 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  registerFile_75 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  registerFile_76 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  registerFile_77 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  registerFile_78 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  registerFile_79 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  registerFile_80 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  registerFile_81 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  registerFile_82 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  registerFile_83 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  registerFile_84 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  registerFile_85 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  registerFile_86 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  registerFile_87 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  registerFile_88 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  registerFile_89 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  registerFile_90 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  registerFile_91 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  registerFile_92 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  registerFile_93 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  registerFile_94 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  registerFile_95 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  registerFile_96 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  registerFile_97 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  registerFile_98 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  registerFile_99 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  registerFile_100 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  registerFile_101 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  registerFile_102 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  registerFile_103 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  registerFile_104 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  registerFile_105 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  registerFile_106 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  registerFile_107 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  registerFile_108 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  registerFile_109 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  registerFile_110 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  registerFile_111 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  registerFile_112 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  registerFile_113 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  registerFile_114 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  registerFile_115 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  registerFile_116 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  registerFile_117 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  registerFile_118 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  registerFile_119 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  registerFile_120 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  registerFile_121 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  registerFile_122 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  registerFile_123 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  registerFile_124 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  registerFile_125 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  registerFile_126 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  registerFile_127 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  registerFile_254 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  registerFile_255 = _RAND_132[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module YM2203(
  input         clock,
  input         reset,
  input         io_cpu_wr,
  input         io_cpu_addr,
  input  [7:0]  io_cpu_din,
  output [7:0]  io_cpu_dout,
  output        io_irq,
  output        io_audio_valid,
  output [15:0] io_audio_bits_psg,
  output [15:0] io_audio_bits_fm
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  m_rst; // @[YM2203.scala 48:17]
  wire  m_clk; // @[YM2203.scala 48:17]
  wire  m_cen; // @[YM2203.scala 48:17]
  wire [7:0] m_din; // @[YM2203.scala 48:17]
  wire  m_addr; // @[YM2203.scala 48:17]
  wire  m_cs_n; // @[YM2203.scala 48:17]
  wire  m_wr_n; // @[YM2203.scala 48:17]
  wire [7:0] m_dout; // @[YM2203.scala 48:17]
  wire  m_irq_n; // @[YM2203.scala 48:17]
  wire [9:0] m_psg_snd; // @[YM2203.scala 48:17]
  wire [15:0] m_fm_snd; // @[YM2203.scala 48:17]
  wire  m_snd_sample; // @[YM2203.scala 48:17]
  reg [15:0] m_io_cen_counter; // @[ClockDivider.scala 40:24]
  wire [16:0] m_io_cen_next = m_io_cen_counter + 16'h2000; // @[ClockDivider.scala 42:19]
  reg  m_io_cen_clockEnable; // @[ClockDivider.scala 41:28]
  jt03 m ( // @[YM2203.scala 48:17]
    .rst(m_rst),
    .clk(m_clk),
    .cen(m_cen),
    .din(m_din),
    .addr(m_addr),
    .cs_n(m_cs_n),
    .wr_n(m_wr_n),
    .dout(m_dout),
    .irq_n(m_irq_n),
    .psg_snd(m_psg_snd),
    .fm_snd(m_fm_snd),
    .snd_sample(m_snd_sample)
  );
  assign io_cpu_dout = m_dout; // @[YM2203.scala 56:15]
  assign io_irq = ~m_irq_n; // @[YM2203.scala 57:13]
  assign io_audio_valid = m_snd_sample; // @[YM2203.scala 58:18]
  assign io_audio_bits_psg = {1'h0,m_psg_snd,5'h0}; // @[YM2203.scala 59:58]
  assign io_audio_bits_fm = m_fm_snd; // @[YM2203.scala 60:20]
  assign m_rst = reset; // @[YM2203.scala 49:21]
  assign m_clk = clock; // @[YM2203.scala 50:21]
  assign m_cen = m_io_cen_clockEnable; // @[YM2203.scala 51:12]
  assign m_din = io_cpu_din; // @[YM2203.scala 55:12]
  assign m_addr = io_cpu_addr; // @[YM2203.scala 54:27]
  assign m_cs_n = 1'h0; // @[YM2203.scala 52:13]
  assign m_wr_n = ~io_cpu_wr; // @[YM2203.scala 53:16]
  always @(posedge clock) begin
    m_io_cen_counter <= m_io_cen_counter + 16'h2000; // @[ClockDivider.scala 40:34]
    m_io_cen_clockEnable <= m_io_cen_next[16]; // @[ClockDivider.scala 41:38]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  m_io_cen_counter = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  m_io_cen_clockEnable = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncReadMemArbiter(
  input         clock,
  input         reset,
  input         io_in_0_rd,
  input  [24:0] io_in_0_addr,
  output [7:0]  io_in_0_dout,
  output        io_in_0_valid,
  input         io_in_1_rd,
  input  [24:0] io_in_1_addr,
  output [7:0]  io_in_1_dout,
  output        io_in_1_wait_n,
  output        io_in_1_valid,
  input         io_in_2_rd,
  input  [24:0] io_in_2_addr,
  output [7:0]  io_in_2_dout,
  input         io_in_3_rd,
  input  [24:0] io_in_3_addr,
  output [7:0]  io_in_3_dout,
  output        io_out_rd,
  output [24:0] io_out_addr,
  input  [7:0]  io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  busyReg; // @[AsyncReadMemArbiter.scala 73:24]
  reg [3:0] indexReg; // @[AsyncReadMemArbiter.scala 74:25]
  wire [3:0] _index_enc_T = io_in_3_rd ? 4'h8 : 4'h0; // @[Mux.scala 47:70]
  wire [3:0] _index_enc_T_1 = io_in_2_rd ? 4'h4 : _index_enc_T; // @[Mux.scala 47:70]
  wire [3:0] _index_enc_T_2 = io_in_1_rd ? 4'h2 : _index_enc_T_1; // @[Mux.scala 47:70]
  wire [3:0] index_enc = io_in_0_rd ? 4'h1 : _index_enc_T_2; // @[Mux.scala 47:70]
  wire [3:0] index = {index_enc[3],index_enc[2],index_enc[1],index_enc[0]}; // @[AsyncReadMemArbiter.scala 77:68]
  wire [3:0] chosen = busyReg ? indexReg : index; // @[AsyncReadMemArbiter.scala 80:19]
  wire  effectiveRequest = ~busyReg & io_out_rd & io_out_wait_n; // @[AsyncReadMemArbiter.scala 83:48]
  wire  _GEN_0 = effectiveRequest | busyReg; // @[AsyncReadMemArbiter.scala 88:32 89:13 73:24]
  wire  io_out_anySelected = chosen[0] | chosen[1] | chosen[2] | chosen[3]; // @[AsyncMemIO.scala 156:45]
  wire [24:0] _io_out_mem_addr_T = chosen[0] ? io_in_0_addr : 25'h0; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_1 = chosen[1] ? io_in_1_addr : 25'h0; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_2 = chosen[2] ? io_in_2_addr : 25'h0; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_3 = chosen[3] ? io_in_3_addr : 25'h0; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_4 = _io_out_mem_addr_T | _io_out_mem_addr_T_1; // @[Mux.scala 27:73]
  wire [24:0] _io_out_mem_addr_T_5 = _io_out_mem_addr_T_4 | _io_out_mem_addr_T_2; // @[Mux.scala 27:73]
  assign io_in_0_dout = io_out_dout; // @[AsyncMemIO.scala 157:19 AsyncReadMemArbiter.scala 96:10]
  assign io_in_0_valid = chosen[0] & io_out_valid; // @[AsyncMemIO.scala 162:30]
  assign io_in_1_dout = io_out_dout; // @[AsyncMemIO.scala 157:19 AsyncReadMemArbiter.scala 96:10]
  assign io_in_1_wait_n = (~io_out_anySelected | chosen[1]) & io_out_wait_n; // @[AsyncMemIO.scala 161:49]
  assign io_in_1_valid = chosen[1] & io_out_valid; // @[AsyncMemIO.scala 162:30]
  assign io_in_2_dout = io_out_dout; // @[AsyncMemIO.scala 157:19 AsyncReadMemArbiter.scala 96:10]
  assign io_in_3_dout = io_out_dout; // @[AsyncMemIO.scala 157:19 AsyncReadMemArbiter.scala 96:10]
  assign io_out_rd = chosen[0] & io_in_0_rd | chosen[1] & io_in_1_rd | chosen[2] & io_in_2_rd | chosen[3] & io_in_3_rd; // @[Mux.scala 27:73]
  assign io_out_addr = _io_out_mem_addr_T_5 | _io_out_mem_addr_T_3; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (reset) begin // @[AsyncReadMemArbiter.scala 73:24]
      busyReg <= 1'h0; // @[AsyncReadMemArbiter.scala 73:24]
    end else if (io_out_valid) begin // @[AsyncReadMemArbiter.scala 86:22]
      busyReg <= 1'h0; // @[AsyncReadMemArbiter.scala 87:13]
    end else begin
      busyReg <= _GEN_0;
    end
    if (reset) begin // @[AsyncReadMemArbiter.scala 74:25]
      indexReg <= 4'h0; // @[AsyncReadMemArbiter.scala 74:25]
    end else if (!(io_out_valid)) begin // @[AsyncReadMemArbiter.scala 86:22]
      if (effectiveRequest) begin // @[AsyncReadMemArbiter.scala 88:32]
        indexReg <= index; // @[AsyncReadMemArbiter.scala 90:14]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busyReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  indexReg = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AudioMixer(
  input         clock,
  input  [13:0] io_in_4,
  input  [13:0] io_in_3,
  input  [15:0] io_in_2,
  input  [15:0] io_in_1,
  input  [15:0] io_in_0,
  output [15:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [21:0] _sum_T_1 = $signed(io_in_0) * 6'sh10; // @[AudioMixer.scala 66:89]
  wire [18:0] _sum_T_3 = $signed(io_in_1) * 3'sh3; // @[AudioMixer.scala 66:89]
  wire [21:0] _sum_T_5 = $signed(io_in_2) * 6'sh10; // @[AudioMixer.scala 66:89]
  wire [15:0] _sum_T_6 = {$signed(io_in_3), 2'h0}; // @[AudioMixer.scala 89:61]
  wire [21:0] _sum_T_7 = $signed(_sum_T_6) * 6'sh1a; // @[AudioMixer.scala 66:89]
  wire [15:0] _sum_T_8 = {$signed(io_in_4), 2'h0}; // @[AudioMixer.scala 89:61]
  wire [21:0] _sum_T_9 = $signed(_sum_T_8) * 6'sh10; // @[AudioMixer.scala 66:89]
  wire [21:0] _GEN_0 = {{3{_sum_T_3[18]}},_sum_T_3}; // @[AudioMixer.scala 67:29]
  wire [22:0] _sum_T_10 = $signed(_sum_T_1) + $signed(_GEN_0); // @[AudioMixer.scala 67:29]
  wire [22:0] _GEN_1 = {{1{_sum_T_5[21]}},_sum_T_5}; // @[AudioMixer.scala 67:29]
  wire [23:0] _sum_T_11 = $signed(_sum_T_10) + $signed(_GEN_1); // @[AudioMixer.scala 67:29]
  wire [23:0] _GEN_2 = {{2{_sum_T_7[21]}},_sum_T_7}; // @[AudioMixer.scala 67:29]
  wire [24:0] _sum_T_12 = $signed(_sum_T_11) + $signed(_GEN_2); // @[AudioMixer.scala 67:29]
  wire [24:0] _GEN_3 = {{3{_sum_T_9[21]}},_sum_T_9}; // @[AudioMixer.scala 67:29]
  wire [25:0] sum = $signed(_sum_T_12) + $signed(_GEN_3); // @[AudioMixer.scala 67:29]
  wire [21:0] io_out_clipped = sum[25:4]; // @[AudioMixer.scala 71:24]
  wire [21:0] _io_out_T_1 = $signed(io_out_clipped) < -22'sh8000 ? $signed(-22'sh8000) : $signed(io_out_clipped); // @[Util.scala 264:51]
  reg [21:0] io_out_REG; // @[AudioMixer.scala 73:12]
  assign io_out = io_out_REG[15:0]; // @[AudioMixer.scala 70:10]
  always @(posedge clock) begin
    if ($signed(_io_out_T_1) < 22'sh7fff) begin // @[Util.scala 264:60]
      if ($signed(io_out_clipped) < -22'sh8000) begin // @[Util.scala 264:51]
        io_out_REG <= -22'sh8000;
      end else begin
        io_out_REG <= io_out_clipped;
      end
    end else begin
      io_out_REG <= 22'sh7fff;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_REG = _RAND_0[21:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Sound(
  input         clock,
  input         reset,
  input         io_ctrl_oki_0_wr,
  input  [15:0] io_ctrl_oki_0_din,
  output [15:0] io_ctrl_oki_0_dout,
  input         io_ctrl_oki_1_wr,
  input  [15:0] io_ctrl_oki_1_din,
  output [15:0] io_ctrl_oki_1_dout,
  input         io_ctrl_nmk_wr,
  input  [22:0] io_ctrl_nmk_addr,
  input  [15:0] io_ctrl_nmk_din,
  input         io_ctrl_ymz_rd,
  input         io_ctrl_ymz_wr,
  input  [22:0] io_ctrl_ymz_addr,
  input  [15:0] io_ctrl_ymz_din,
  output [15:0] io_ctrl_ymz_dout,
  input         io_ctrl_req,
  input  [15:0] io_ctrl_data,
  output        io_ctrl_irq,
  input  [3:0]  io_gameIndex,
  input  [1:0]  io_gameConfig_sound_0_device,
  output        io_rom_0_rd,
  output [24:0] io_rom_0_addr,
  input  [7:0]  io_rom_0_dout,
  input         io_rom_0_wait_n,
  input         io_rom_0_valid,
  output [24:0] io_rom_1_addr,
  input  [7:0]  io_rom_1_dout,
  input         io_rom_1_valid,
  output [15:0] io_audio
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  cpu_clock; // @[Sound.scala 74:19]
  wire  cpu_reset; // @[Sound.scala 74:19]
  wire [15:0] cpu_io_addr; // @[Sound.scala 74:19]
  wire [7:0] cpu_io_din; // @[Sound.scala 74:19]
  wire [7:0] cpu_io_dout; // @[Sound.scala 74:19]
  wire  cpu_io_rd; // @[Sound.scala 74:19]
  wire  cpu_io_wr; // @[Sound.scala 74:19]
  wire  cpu_io_rfsh; // @[Sound.scala 74:19]
  wire  cpu_io_mreq; // @[Sound.scala 74:19]
  wire  cpu_io_iorq; // @[Sound.scala 74:19]
  wire  cpu_io_int; // @[Sound.scala 74:19]
  wire  cpu_io_nmi; // @[Sound.scala 74:19]
  wire  soundRam_clock; // @[Sound.scala 83:24]
  wire  soundRam_io_rd; // @[Sound.scala 83:24]
  wire  soundRam_io_wr; // @[Sound.scala 83:24]
  wire [12:0] soundRam_io_addr; // @[Sound.scala 83:24]
  wire [7:0] soundRam_io_din; // @[Sound.scala 83:24]
  wire [7:0] soundRam_io_dout; // @[Sound.scala 83:24]
  wire  nmk_clock; // @[Sound.scala 90:19]
  wire  nmk_io_cpu_wr; // @[Sound.scala 90:19]
  wire [22:0] nmk_io_cpu_addr; // @[Sound.scala 90:19]
  wire [15:0] nmk_io_cpu_din; // @[Sound.scala 90:19]
  wire [24:0] nmk_io_addr_0_in; // @[Sound.scala 90:19]
  wire [24:0] nmk_io_addr_0_out; // @[Sound.scala 90:19]
  wire [24:0] nmk_io_addr_1_in; // @[Sound.scala 90:19]
  wire [24:0] nmk_io_addr_1_out; // @[Sound.scala 90:19]
  wire  oki_0_clock; // @[Sound.scala 96:21]
  wire  oki_0_reset; // @[Sound.scala 96:21]
  wire  oki_0_io_cpu_wr; // @[Sound.scala 96:21]
  wire [7:0] oki_0_io_cpu_din; // @[Sound.scala 96:21]
  wire [7:0] oki_0_io_cpu_dout; // @[Sound.scala 96:21]
  wire [17:0] oki_0_io_rom_addr; // @[Sound.scala 96:21]
  wire [7:0] oki_0_io_rom_dout; // @[Sound.scala 96:21]
  wire  oki_0_io_rom_valid; // @[Sound.scala 96:21]
  wire  oki_0_io_audio_valid; // @[Sound.scala 96:21]
  wire [13:0] oki_0_io_audio_bits; // @[Sound.scala 96:21]
  wire  oki_1_clock; // @[Sound.scala 96:21]
  wire  oki_1_reset; // @[Sound.scala 96:21]
  wire  oki_1_io_cpu_wr; // @[Sound.scala 96:21]
  wire [7:0] oki_1_io_cpu_din; // @[Sound.scala 96:21]
  wire [7:0] oki_1_io_cpu_dout; // @[Sound.scala 96:21]
  wire [17:0] oki_1_io_rom_addr; // @[Sound.scala 96:21]
  wire [7:0] oki_1_io_rom_dout; // @[Sound.scala 96:21]
  wire  oki_1_io_rom_valid; // @[Sound.scala 96:21]
  wire  oki_1_io_audio_valid; // @[Sound.scala 96:21]
  wire [13:0] oki_1_io_audio_bits; // @[Sound.scala 96:21]
  wire  ymz280b_clock; // @[Sound.scala 102:23]
  wire  ymz280b_reset; // @[Sound.scala 102:23]
  wire  ymz280b_io_cpu_rd; // @[Sound.scala 102:23]
  wire  ymz280b_io_cpu_wr; // @[Sound.scala 102:23]
  wire  ymz280b_io_cpu_addr; // @[Sound.scala 102:23]
  wire [7:0] ymz280b_io_cpu_din; // @[Sound.scala 102:23]
  wire [7:0] ymz280b_io_cpu_dout; // @[Sound.scala 102:23]
  wire  ymz280b_io_rom_rd; // @[Sound.scala 102:23]
  wire [23:0] ymz280b_io_rom_addr; // @[Sound.scala 102:23]
  wire [7:0] ymz280b_io_rom_dout; // @[Sound.scala 102:23]
  wire  ymz280b_io_rom_wait_n; // @[Sound.scala 102:23]
  wire  ymz280b_io_rom_valid; // @[Sound.scala 102:23]
  wire  ymz280b_io_audio_valid; // @[Sound.scala 102:23]
  wire [15:0] ymz280b_io_audio_bits_left; // @[Sound.scala 102:23]
  wire  ymz280b_io_irq; // @[Sound.scala 102:23]
  wire  ym2203_clock; // @[Sound.scala 108:22]
  wire  ym2203_reset; // @[Sound.scala 108:22]
  wire  ym2203_io_cpu_wr; // @[Sound.scala 108:22]
  wire  ym2203_io_cpu_addr; // @[Sound.scala 108:22]
  wire [7:0] ym2203_io_cpu_din; // @[Sound.scala 108:22]
  wire [7:0] ym2203_io_cpu_dout; // @[Sound.scala 108:22]
  wire  ym2203_io_irq; // @[Sound.scala 108:22]
  wire  ym2203_io_audio_valid; // @[Sound.scala 108:22]
  wire [15:0] ym2203_io_audio_bits_psg; // @[Sound.scala 108:22]
  wire [15:0] ym2203_io_audio_bits_fm; // @[Sound.scala 108:22]
  wire  arbiter_clock; // @[Sound.scala 119:23]
  wire  arbiter_reset; // @[Sound.scala 119:23]
  wire  arbiter_io_in_0_rd; // @[Sound.scala 119:23]
  wire [24:0] arbiter_io_in_0_addr; // @[Sound.scala 119:23]
  wire [7:0] arbiter_io_in_0_dout; // @[Sound.scala 119:23]
  wire  arbiter_io_in_0_valid; // @[Sound.scala 119:23]
  wire  arbiter_io_in_1_rd; // @[Sound.scala 119:23]
  wire [24:0] arbiter_io_in_1_addr; // @[Sound.scala 119:23]
  wire [7:0] arbiter_io_in_1_dout; // @[Sound.scala 119:23]
  wire  arbiter_io_in_1_wait_n; // @[Sound.scala 119:23]
  wire  arbiter_io_in_1_valid; // @[Sound.scala 119:23]
  wire  arbiter_io_in_2_rd; // @[Sound.scala 119:23]
  wire [24:0] arbiter_io_in_2_addr; // @[Sound.scala 119:23]
  wire [7:0] arbiter_io_in_2_dout; // @[Sound.scala 119:23]
  wire  arbiter_io_in_3_rd; // @[Sound.scala 119:23]
  wire [24:0] arbiter_io_in_3_addr; // @[Sound.scala 119:23]
  wire [7:0] arbiter_io_in_3_dout; // @[Sound.scala 119:23]
  wire  arbiter_io_out_rd; // @[Sound.scala 119:23]
  wire [24:0] arbiter_io_out_addr; // @[Sound.scala 119:23]
  wire [7:0] arbiter_io_out_dout; // @[Sound.scala 119:23]
  wire  arbiter_io_out_wait_n; // @[Sound.scala 119:23]
  wire  arbiter_io_out_valid; // @[Sound.scala 119:23]
  wire  io_audio_mixer_clock; // @[AudioMixer.scala 100:23]
  wire [13:0] io_audio_mixer_io_in_4; // @[AudioMixer.scala 100:23]
  wire [13:0] io_audio_mixer_io_in_3; // @[AudioMixer.scala 100:23]
  wire [15:0] io_audio_mixer_io_in_2; // @[AudioMixer.scala 100:23]
  wire [15:0] io_audio_mixer_io_in_1; // @[AudioMixer.scala 100:23]
  wire [15:0] io_audio_mixer_io_in_0; // @[AudioMixer.scala 100:23]
  wire [15:0] io_audio_mixer_io_out; // @[AudioMixer.scala 100:23]
  reg  reqReg; // @[Reg.scala 35:20]
  wire  _GEN_0 = io_ctrl_req | reqReg; // @[Reg.scala 36:18 35:20 36:22]
  reg [15:0] dataReg; // @[Reg.scala 19:16]
  reg [3:0] z80BankReg; // @[Sound.scala 69:27]
  reg [3:0] okiBankHiReg; // @[Sound.scala 70:29]
  reg [3:0] okiBankLoReg; // @[Sound.scala 71:29]
  wire [3:0] mem_bank = oki_0_io_rom_addr[17] ? okiBankHiReg : okiBankLoReg; // @[Sound.scala 146:19]
  wire [20:0] _mem_T_2 = {mem_bank,oki_0_io_rom_addr[16:0]}; // @[Sound.scala 149:12]
  wire  _T_1 = io_gameConfig_sound_0_device == 2'h1; // @[Sound.scala 122:57]
  wire  _T_2 = io_gameConfig_sound_0_device == 2'h3; // @[Sound.scala 123:50]
  wire [15:0] addr = cpu_io_addr; // @[MemMap.scala 76:25]
  wire  cs = addr <= 16'h3fff; // @[Util.scala 64:72]
  wire  _progRom_rd_T = ~cpu_io_rfsh; // @[MemMap.scala 117:23]
  wire  progRom_rd = io_gameIndex == 4'h7 & (cs & ~cpu_io_rfsh); // @[MemMap.scala 117:14 Sound.scala 165:42 MemIO.scala 83:8]
  wire  cs_1 = addr >= 16'h4000 & addr <= 16'h7fff; // @[Util.scala 64:67]
  wire  bankRom_rd = io_gameIndex == 4'h7 & (cs_1 & ~cpu_io_rfsh); // @[MemMap.scala 117:14 Sound.scala 165:42 MemIO.scala 83:8]
  wire [3:0] mem_bank_1 = oki_1_io_rom_addr[17] ? okiBankHiReg : okiBankLoReg; // @[Sound.scala 146:19]
  wire [20:0] _mem_T_6 = {mem_bank_1,oki_1_io_rom_addr[16:0]}; // @[Sound.scala 149:12]
  wire [7:0] mem_3_dout = arbiter_io_in_2_dout; // @[AsyncMemIO.scala 134:19 AsyncReadMemArbiter.scala 68:54]
  wire [17:0] _bankRom_addr_T_1 = {z80BankReg,addr[13:0]}; // @[Sound.scala 167:69]
  wire [7:0] mem_4_dout = arbiter_io_in_3_dout; // @[AsyncMemIO.scala 134:19 AsyncReadMemArbiter.scala 68:54]
  wire [7:0] _GEN_3 = cs_1 & cpu_io_mreq & cpu_io_rd ? mem_4_dout : mem_3_dout; // @[MemMap.scala 119:{38,48}]
  wire  cs_2 = addr >= 16'he000; // @[Util.scala 64:58]
  wire  _soundRam_io_wr_T = cs_2 & cpu_io_mreq; // @[MemMap.scala 97:20]
  wire [7:0] _GEN_4 = _soundRam_io_wr_T & cpu_io_rd ? soundRam_io_dout : _GEN_3; // @[MemMap.scala 100:{38,48}]
  wire [15:0] addr_3 = cpu_io_addr & 16'hff; // @[IOMap.scala 76:25]
  wire  cs_3 = addr_3 <= 16'h0; // @[Util.scala 64:72]
  wire  cs_4 = addr_3 >= 16'h30 & addr_3 <= 16'h30; // @[Util.scala 64:67]
  wire [7:0] _GEN_7 = cs_4 & cpu_io_iorq & cpu_io_rd ? dataReg[7:0] : _GEN_4; // @[IOMap.scala 163:{38,48}]
  wire  cs_5 = addr_3 >= 16'h40 & addr_3 <= 16'h40; // @[Util.scala 64:67]
  wire [7:0] _GEN_9 = cs_5 & cpu_io_iorq & cpu_io_rd ? dataReg[15:8] : _GEN_7; // @[IOMap.scala 163:{38,48}]
  wire  cs_6 = addr_3 >= 16'h50 & addr_3 <= 16'h51; // @[Util.scala 64:67]
  wire  _ym2203_io_cpu_wr_T = cs_6 & cpu_io_iorq; // @[IOMap.scala 97:20]
  wire [7:0] _GEN_10 = _ym2203_io_cpu_wr_T & cpu_io_rd ? ym2203_io_cpu_dout : _GEN_9; // @[IOMap.scala 100:{38,48}]
  wire  cs_7 = addr_3 >= 16'h60 & addr_3 <= 16'h60; // @[Util.scala 64:67]
  wire  _oki_1_io_cpu_wr_T = cs_7 & cpu_io_iorq; // @[IOMap.scala 97:20]
  wire  cs_8 = addr_3 >= 16'h70 & addr_3 <= 16'h70; // @[Util.scala 64:67]
  wire [3:0] _okiBankHiReg_T_1 = cpu_io_dout[7:4] & 4'h3; // @[Sound.scala 160:32]
  wire [3:0] _okiBankLoReg_T_1 = cpu_io_dout[3:0] & 4'h3; // @[Sound.scala 161:32]
  wire [15:0] _GEN_31 = io_gameIndex == 4'h7 ? {{8'd0}, cpu_io_dout} : io_ctrl_oki_1_din; // @[Sound.scala 165:42 IOMap.scala 99:15 Sound.scala 97:16]
  reg [15:0] io_audio_r; // @[Reg.scala 19:16]
  reg [15:0] io_audio_r_1; // @[Reg.scala 19:16]
  reg [15:0] io_audio_r_2; // @[Reg.scala 19:16]
  reg [13:0] io_audio_r_3; // @[Reg.scala 19:16]
  reg [13:0] io_audio_r_4; // @[Reg.scala 19:16]
  wire [23:0] mem_2_addr = ymz280b_io_rom_addr; // @[AsyncMemIO.scala 134:19 138:14]
  CPU_1 cpu ( // @[Sound.scala 74:19]
    .clock(cpu_clock),
    .reset(cpu_reset),
    .io_addr(cpu_io_addr),
    .io_din(cpu_io_din),
    .io_dout(cpu_io_dout),
    .io_rd(cpu_io_rd),
    .io_wr(cpu_io_wr),
    .io_rfsh(cpu_io_rfsh),
    .io_mreq(cpu_io_mreq),
    .io_iorq(cpu_io_iorq),
    .io_int(cpu_io_int),
    .io_nmi(cpu_io_nmi)
  );
  SinglePortRam_1 soundRam ( // @[Sound.scala 83:24]
    .clock(soundRam_clock),
    .io_rd(soundRam_io_rd),
    .io_wr(soundRam_io_wr),
    .io_addr(soundRam_io_addr),
    .io_din(soundRam_io_din),
    .io_dout(soundRam_io_dout)
  );
  NMK112 nmk ( // @[Sound.scala 90:19]
    .clock(nmk_clock),
    .io_cpu_wr(nmk_io_cpu_wr),
    .io_cpu_addr(nmk_io_cpu_addr),
    .io_cpu_din(nmk_io_cpu_din),
    .io_addr_0_in(nmk_io_addr_0_in),
    .io_addr_0_out(nmk_io_addr_0_out),
    .io_addr_1_in(nmk_io_addr_1_in),
    .io_addr_1_out(nmk_io_addr_1_out)
  );
  OKIM6295 oki_0 ( // @[Sound.scala 96:21]
    .clock(oki_0_clock),
    .reset(oki_0_reset),
    .io_cpu_wr(oki_0_io_cpu_wr),
    .io_cpu_din(oki_0_io_cpu_din),
    .io_cpu_dout(oki_0_io_cpu_dout),
    .io_rom_addr(oki_0_io_rom_addr),
    .io_rom_dout(oki_0_io_rom_dout),
    .io_rom_valid(oki_0_io_rom_valid),
    .io_audio_valid(oki_0_io_audio_valid),
    .io_audio_bits(oki_0_io_audio_bits)
  );
  OKIM6295_1 oki_1 ( // @[Sound.scala 96:21]
    .clock(oki_1_clock),
    .reset(oki_1_reset),
    .io_cpu_wr(oki_1_io_cpu_wr),
    .io_cpu_din(oki_1_io_cpu_din),
    .io_cpu_dout(oki_1_io_cpu_dout),
    .io_rom_addr(oki_1_io_rom_addr),
    .io_rom_dout(oki_1_io_rom_dout),
    .io_rom_valid(oki_1_io_rom_valid),
    .io_audio_valid(oki_1_io_audio_valid),
    .io_audio_bits(oki_1_io_audio_bits)
  );
  YMZ280B ymz280b ( // @[Sound.scala 102:23]
    .clock(ymz280b_clock),
    .reset(ymz280b_reset),
    .io_cpu_rd(ymz280b_io_cpu_rd),
    .io_cpu_wr(ymz280b_io_cpu_wr),
    .io_cpu_addr(ymz280b_io_cpu_addr),
    .io_cpu_din(ymz280b_io_cpu_din),
    .io_cpu_dout(ymz280b_io_cpu_dout),
    .io_rom_rd(ymz280b_io_rom_rd),
    .io_rom_addr(ymz280b_io_rom_addr),
    .io_rom_dout(ymz280b_io_rom_dout),
    .io_rom_wait_n(ymz280b_io_rom_wait_n),
    .io_rom_valid(ymz280b_io_rom_valid),
    .io_audio_valid(ymz280b_io_audio_valid),
    .io_audio_bits_left(ymz280b_io_audio_bits_left),
    .io_irq(ymz280b_io_irq)
  );
  YM2203 ym2203 ( // @[Sound.scala 108:22]
    .clock(ym2203_clock),
    .reset(ym2203_reset),
    .io_cpu_wr(ym2203_io_cpu_wr),
    .io_cpu_addr(ym2203_io_cpu_addr),
    .io_cpu_din(ym2203_io_cpu_din),
    .io_cpu_dout(ym2203_io_cpu_dout),
    .io_irq(ym2203_io_irq),
    .io_audio_valid(ym2203_io_audio_valid),
    .io_audio_bits_psg(ym2203_io_audio_bits_psg),
    .io_audio_bits_fm(ym2203_io_audio_bits_fm)
  );
  AsyncReadMemArbiter arbiter ( // @[Sound.scala 119:23]
    .clock(arbiter_clock),
    .reset(arbiter_reset),
    .io_in_0_rd(arbiter_io_in_0_rd),
    .io_in_0_addr(arbiter_io_in_0_addr),
    .io_in_0_dout(arbiter_io_in_0_dout),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_1_rd(arbiter_io_in_1_rd),
    .io_in_1_addr(arbiter_io_in_1_addr),
    .io_in_1_dout(arbiter_io_in_1_dout),
    .io_in_1_wait_n(arbiter_io_in_1_wait_n),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_2_rd(arbiter_io_in_2_rd),
    .io_in_2_addr(arbiter_io_in_2_addr),
    .io_in_2_dout(arbiter_io_in_2_dout),
    .io_in_3_rd(arbiter_io_in_3_rd),
    .io_in_3_addr(arbiter_io_in_3_addr),
    .io_in_3_dout(arbiter_io_in_3_dout),
    .io_out_rd(arbiter_io_out_rd),
    .io_out_addr(arbiter_io_out_addr),
    .io_out_dout(arbiter_io_out_dout),
    .io_out_wait_n(arbiter_io_out_wait_n),
    .io_out_valid(arbiter_io_out_valid)
  );
  AudioMixer io_audio_mixer ( // @[AudioMixer.scala 100:23]
    .clock(io_audio_mixer_clock),
    .io_in_4(io_audio_mixer_io_in_4),
    .io_in_3(io_audio_mixer_io_in_3),
    .io_in_2(io_audio_mixer_io_in_2),
    .io_in_1(io_audio_mixer_io_in_1),
    .io_in_0(io_audio_mixer_io_in_0),
    .io_out(io_audio_mixer_io_out)
  );
  assign io_ctrl_oki_0_dout = {{8'd0}, oki_0_io_cpu_dout}; // @[Sound.scala 97:16]
  assign io_ctrl_oki_1_dout = {{8'd0}, oki_1_io_cpu_dout}; // @[Sound.scala 97:16]
  assign io_ctrl_ymz_dout = {{8'd0}, ymz280b_io_cpu_dout}; // @[Sound.scala 103:18]
  assign io_ctrl_irq = ymz280b_io_irq; // @[Sound.scala 105:15]
  assign io_rom_0_rd = arbiter_io_out_rd; // @[Sound.scala 125:5]
  assign io_rom_0_addr = arbiter_io_out_addr; // @[Sound.scala 125:5]
  assign io_rom_1_addr = io_gameIndex == 4'h2 ? nmk_io_addr_1_out : {{4'd0}, _mem_T_6}; // @[Sound.scala 147:8]
  assign io_audio = io_audio_mixer_io_out; // @[Sound.scala 179:12]
  assign cpu_clock = clock;
  assign cpu_reset = reset;
  assign cpu_io_din = _oki_1_io_cpu_wr_T & cpu_io_rd ? oki_1_io_cpu_dout : _GEN_10; // @[IOMap.scala 100:{38,48}]
  assign cpu_io_int = ym2203_io_irq; // @[Sound.scala 64:17 109:7]
  assign cpu_io_nmi = reqReg; // @[Sound.scala 80:14]
  assign soundRam_clock = clock;
  assign soundRam_io_rd = io_gameIndex == 4'h7 & (cs_2 & _progRom_rd_T); // @[Sound.scala 165:42 MemMap.scala 96:14 MemIO.scala 317:8]
  assign soundRam_io_wr = io_gameIndex == 4'h7 & (cs_2 & cpu_io_mreq & cpu_io_wr); // @[Sound.scala 165:42 MemMap.scala 97:14 MemIO.scala 318:8]
  assign soundRam_io_addr = addr[12:0];
  assign soundRam_io_din = cpu_io_dout; // @[Sound.scala 165:42 MemMap.scala 99:15]
  assign nmk_clock = clock;
  assign nmk_io_cpu_wr = io_ctrl_nmk_wr; // @[Sound.scala 91:14]
  assign nmk_io_cpu_addr = io_ctrl_nmk_addr; // @[Sound.scala 91:14]
  assign nmk_io_cpu_din = io_ctrl_nmk_din; // @[Sound.scala 91:14]
  assign nmk_io_addr_0_in = {{7'd0}, oki_0_io_rom_addr}; // @[NMK112.scala 80:22]
  assign nmk_io_addr_1_in = {{7'd0}, oki_1_io_rom_addr}; // @[NMK112.scala 80:22]
  assign oki_0_clock = clock;
  assign oki_0_reset = reset;
  assign oki_0_io_cpu_wr = io_ctrl_oki_0_wr; // @[Sound.scala 97:16]
  assign oki_0_io_cpu_din = io_ctrl_oki_0_din[7:0]; // @[Sound.scala 97:16]
  assign oki_0_io_rom_dout = arbiter_io_in_0_dout; // @[AsyncMemIO.scala 134:19 AsyncReadMemArbiter.scala 68:54]
  assign oki_0_io_rom_valid = arbiter_io_in_0_valid; // @[AsyncMemIO.scala 134:19 AsyncReadMemArbiter.scala 68:54]
  assign oki_1_clock = clock;
  assign oki_1_reset = reset;
  assign oki_1_io_cpu_wr = io_gameIndex == 4'h7 ? cs_7 & cpu_io_iorq & cpu_io_wr : io_ctrl_oki_1_wr; // @[Sound.scala 165:42 IOMap.scala 97:14 Sound.scala 97:16]
  assign oki_1_io_cpu_din = _GEN_31[7:0];
  assign oki_1_io_rom_dout = io_rom_1_dout; // @[AsyncMemIO.scala 104:19 Sound.scala 128:40]
  assign oki_1_io_rom_valid = io_rom_1_valid; // @[AsyncMemIO.scala 104:19 Sound.scala 128:40]
  assign ymz280b_clock = clock;
  assign ymz280b_reset = reset;
  assign ymz280b_io_cpu_rd = io_ctrl_ymz_rd; // @[Sound.scala 103:18]
  assign ymz280b_io_cpu_wr = io_ctrl_ymz_wr; // @[Sound.scala 103:18]
  assign ymz280b_io_cpu_addr = io_ctrl_ymz_addr[0]; // @[Sound.scala 103:18]
  assign ymz280b_io_cpu_din = io_ctrl_ymz_din[7:0]; // @[Sound.scala 103:18]
  assign ymz280b_io_rom_dout = arbiter_io_in_1_dout; // @[AsyncMemIO.scala 134:19 AsyncReadMemArbiter.scala 68:54]
  assign ymz280b_io_rom_wait_n = arbiter_io_in_1_wait_n; // @[AsyncMemIO.scala 134:19 AsyncReadMemArbiter.scala 68:54]
  assign ymz280b_io_rom_valid = arbiter_io_in_1_valid; // @[AsyncMemIO.scala 134:19 AsyncReadMemArbiter.scala 68:54]
  assign ym2203_clock = clock;
  assign ym2203_reset = reset;
  assign ym2203_io_cpu_wr = io_gameIndex == 4'h7 & (cs_6 & cpu_io_iorq & cpu_io_wr); // @[Sound.scala 165:42 IOMap.scala 97:14 MemIO.scala 318:8]
  assign ym2203_io_cpu_addr = addr_3[0];
  assign ym2203_io_cpu_din = cpu_io_dout; // @[Sound.scala 165:42 MemMap.scala 99:15]
  assign arbiter_clock = clock;
  assign arbiter_reset = reset;
  assign arbiter_io_in_0_rd = io_gameConfig_sound_0_device == 2'h2; // @[Sound.scala 121:79]
  assign arbiter_io_in_0_addr = io_gameIndex == 4'h2 ? nmk_io_addr_0_out : {{4'd0}, _mem_T_2}; // @[Sound.scala 147:8]
  assign arbiter_io_in_1_rd = _T_1 & ymz280b_io_rom_rd; // @[AsyncMemIO.scala 135:21]
  assign arbiter_io_in_1_addr = {{1'd0}, mem_2_addr}; // @[AsyncReadMemArbiter.scala 68:54]
  assign arbiter_io_in_2_rd = _T_2 & progRom_rd; // @[AsyncMemIO.scala 135:21]
  assign arbiter_io_in_2_addr = {{9'd0}, addr}; // @[Sound.scala 113:21]
  assign arbiter_io_in_3_rd = _T_2 & bankRom_rd; // @[AsyncMemIO.scala 135:21]
  assign arbiter_io_in_3_addr = {{7'd0}, _bankRom_addr_T_1}; // @[Sound.scala 114:21]
  assign arbiter_io_out_dout = io_rom_0_dout; // @[Sound.scala 125:5]
  assign arbiter_io_out_wait_n = io_rom_0_wait_n; // @[Sound.scala 125:5]
  assign arbiter_io_out_valid = io_rom_0_valid; // @[Sound.scala 125:5]
  assign io_audio_mixer_clock = clock;
  assign io_audio_mixer_io_in_4 = io_audio_r_4; // @[MixedVec.scala 117:9]
  assign io_audio_mixer_io_in_3 = io_audio_r_3; // @[MixedVec.scala 117:9]
  assign io_audio_mixer_io_in_2 = io_audio_r_2; // @[MixedVec.scala 117:9]
  assign io_audio_mixer_io_in_1 = io_audio_r_1; // @[MixedVec.scala 117:9]
  assign io_audio_mixer_io_in_0 = io_audio_r; // @[MixedVec.scala 117:9]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      reqReg <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_gameIndex == 4'h7) begin // @[Sound.scala 165:42]
      if (cs_5 & cpu_io_iorq & cpu_io_rd) begin // @[IOMap.scala 163:38]
        reqReg <= 1'h0; // @[Sound.scala 136:12]
      end else if (cs_4 & cpu_io_iorq & cpu_io_rd) begin // @[IOMap.scala 163:38]
        reqReg <= 1'h0; // @[Sound.scala 136:12]
      end else begin
        reqReg <= _GEN_0;
      end
    end else begin
      reqReg <= _GEN_0;
    end
    if (io_ctrl_req) begin // @[Reg.scala 20:18]
      dataReg <= io_ctrl_data; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[Sound.scala 69:27]
      z80BankReg <= 4'h0; // @[Sound.scala 69:27]
    end else if (io_gameIndex == 4'h7) begin // @[Sound.scala 165:42]
      if (cs_3 & cpu_io_iorq & cpu_io_wr) begin // @[IOMap.scala 172:38]
        z80BankReg <= cpu_io_dout[3:0]; // @[Sound.scala 170:48]
      end
    end
    if (reset) begin // @[Sound.scala 70:29]
      okiBankHiReg <= 4'h0; // @[Sound.scala 70:29]
    end else if (io_gameIndex == 4'h7) begin // @[Sound.scala 165:42]
      if (cs_8 & cpu_io_iorq & cpu_io_wr) begin // @[IOMap.scala 172:38]
        okiBankHiReg <= _okiBankHiReg_T_1; // @[Sound.scala 160:18]
      end
    end
    if (reset) begin // @[Sound.scala 71:29]
      okiBankLoReg <= 4'h0; // @[Sound.scala 71:29]
    end else if (io_gameIndex == 4'h7) begin // @[Sound.scala 165:42]
      if (cs_8 & cpu_io_iorq & cpu_io_wr) begin // @[IOMap.scala 172:38]
        okiBankLoReg <= _okiBankLoReg_T_1; // @[Sound.scala 161:18]
      end
    end
    if (ymz280b_io_audio_valid) begin // @[Reg.scala 20:18]
      io_audio_r <= ymz280b_io_audio_bits_left; // @[Reg.scala 20:22]
    end
    if (ym2203_io_audio_valid) begin // @[Reg.scala 20:18]
      io_audio_r_1 <= ym2203_io_audio_bits_psg; // @[Reg.scala 20:22]
    end
    if (ym2203_io_audio_valid) begin // @[Reg.scala 20:18]
      io_audio_r_2 <= ym2203_io_audio_bits_fm; // @[Reg.scala 20:22]
    end
    if (oki_0_io_audio_valid) begin // @[Reg.scala 20:18]
      io_audio_r_3 <= oki_0_io_audio_bits; // @[Reg.scala 20:22]
    end
    if (oki_1_io_audio_valid) begin // @[Reg.scala 20:18]
      io_audio_r_4 <= oki_1_io_audio_bits; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reqReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  dataReg = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  z80BankReg = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  okiBankHiReg = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  okiBankLoReg = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  io_audio_r = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  io_audio_r_1 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  io_audio_r_2 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  io_audio_r_3 = _RAND_8[13:0];
  _RAND_9 = {1{`RANDOM}};
  io_audio_r_4 = _RAND_9[13:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReadDataFreezer_1(
  input         clock,
  input         reset,
  input         io_targetClock,
  input         io_in_rd,
  input  [24:0] io_in_addr,
  output [7:0]  io_in_dout,
  output        io_in_wait_n,
  output        io_in_valid,
  output        io_out_rd,
  output [24:0] io_out_addr,
  input  [7:0]  io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  clear_s; // @[Util.scala 242:26]
  wire  _clear_s_dataReg_T = ~clear_s; // @[Util.scala 243:31]
  reg  clear_REG; // @[Util.scala 151:40]
  wire  clear = clear_s ^ clear_REG; // @[Util.scala 151:31]
  reg  wait_n_enableReg; // @[Util.scala 188:28]
  wire  _GEN_1 = clear ? 1'h0 : wait_n_enableReg; // @[Util.scala 188:28 189:{53,65}]
  wire  _GEN_2 = io_out_wait_n | _GEN_1; // @[Util.scala 189:{13,25}]
  wire  _wait_n_T = ~clear; // @[Util.scala 190:24]
  reg  valid_enableReg; // @[Util.scala 188:28]
  wire  _GEN_3 = clear ? 1'h0 : valid_enableReg; // @[Util.scala 188:28 189:{53,65}]
  wire  _GEN_4 = io_out_valid | _GEN_3; // @[Util.scala 189:{13,25}]
  reg [7:0] data_dataReg; // @[Reg.scala 19:16]
  reg  data_enableReg; // @[Util.scala 204:28]
  wire  _GEN_6 = io_out_valid | data_enableReg; // @[Util.scala 204:28 205:{54,66}]
  reg  pendingRead; // @[Crossing.scala 116:28]
  wire  effectiveRead = io_in_rd & io_out_wait_n; // @[Crossing.scala 117:32]
  reg  clearRead_REG; // @[Crossing.scala 118:35]
  wire  clearRead = clear & clearRead_REG; // @[Crossing.scala 118:25]
  wire  _GEN_8 = clearRead ? 1'h0 : pendingRead; // @[Crossing.scala 116:28 119:{69,83}]
  wire  _GEN_9 = effectiveRead | _GEN_8; // @[Crossing.scala 119:{23,37}]
  assign io_in_dout = data_enableReg & _wait_n_T ? data_dataReg : io_out_dout; // @[Util.scala 206:8]
  assign io_in_wait_n = io_out_wait_n | wait_n_enableReg & ~clear; // @[Util.scala 190:7]
  assign io_in_valid = io_out_valid | valid_enableReg & ~clear; // @[Util.scala 190:7]
  assign io_out_rd = io_in_rd & (~pendingRead | clearRead); // @[Crossing.scala 128:25]
  assign io_out_addr = io_in_addr; // @[Crossing.scala 122:9]
  always @(posedge io_targetClock) begin
    if (reset) begin // @[Util.scala 242:26]
      clear_s <= 1'h0; // @[Util.scala 242:26]
    end else begin
      clear_s <= _clear_s_dataReg_T;
    end
  end
  always @(posedge clock) begin
    clear_REG <= clear_s; // @[Util.scala 151:40]
    if (reset) begin // @[Util.scala 188:28]
      wait_n_enableReg <= 1'h0; // @[Util.scala 188:28]
    end else begin
      wait_n_enableReg <= _GEN_2;
    end
    if (reset) begin // @[Util.scala 188:28]
      valid_enableReg <= 1'h0; // @[Util.scala 188:28]
    end else begin
      valid_enableReg <= _GEN_4;
    end
    if (io_out_valid) begin // @[Reg.scala 20:18]
      data_dataReg <= io_out_dout; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[Util.scala 204:28]
      data_enableReg <= 1'h0; // @[Util.scala 204:28]
    end else if (clear) begin // @[Util.scala 205:17]
      data_enableReg <= 1'h0; // @[Util.scala 205:29]
    end else begin
      data_enableReg <= _GEN_6;
    end
    if (reset) begin // @[Crossing.scala 116:28]
      pendingRead <= 1'h0; // @[Crossing.scala 116:28]
    end else begin
      pendingRead <= _GEN_9;
    end
    clearRead_REG <= io_out_valid | valid_enableReg & ~clear; // @[Util.scala 190:7]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  clear_s = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  clear_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wait_n_enableReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  valid_enableReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  data_dataReg = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_enableReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pendingRead = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  clearRead_REG = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits,
  output [6:0]  io_count,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:63]; // @[Decoupled.scala 275:44]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:44]
  wire [5:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:44]
  wire [63:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:44]
  wire [63:0] ram_MPORT_data; // @[Decoupled.scala 275:44]
  wire [5:0] ram_MPORT_addr; // @[Decoupled.scala 275:44]
  wire  ram_MPORT_mask; // @[Decoupled.scala 275:44]
  wire  ram_MPORT_en; // @[Decoupled.scala 275:44]
  reg  ram_io_deq_bits_MPORT_en_pipe_0;
  reg [5:0] ram_io_deq_bits_MPORT_addr_pipe_0;
  reg [5:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [5:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 278:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 279:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 280:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 281:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  wire [5:0] _value_T_1 = enq_ptr_value + 6'h1; // @[Counter.scala 77:24]
  wire [5:0] _value_T_3 = deq_ptr_value + 6'h1; // @[Counter.scala 77:24]
  wire [6:0] _deq_ptr_next_T_1 = 7'h40 - 7'h1; // @[Decoupled.scala 308:57]
  wire [6:0] _GEN_15 = {{1'd0}, deq_ptr_value}; // @[Decoupled.scala 308:42]
  wire [5:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 328:32]
  wire [6:0] _io_count_T_1 = maybe_full & ptr_match ? 7'h40 : 7'h0; // @[Decoupled.scala 331:20]
  wire [6:0] _GEN_16 = {{1'd0}, ptr_diff}; // @[Decoupled.scala 331:62]
  assign ram_io_deq_bits_MPORT_en = ram_io_deq_bits_MPORT_en_pipe_0;
  assign ram_io_deq_bits_MPORT_addr = ram_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:44]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 305:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 304:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_count = _io_count_T_1 | _GEN_16; // @[Decoupled.scala 331:62]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 275:44]
    end
    ram_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_15 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 308:27]
          ram_io_deq_bits_MPORT_addr_pipe_0 <= 6'h0;
        end else begin
          ram_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 6'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 298:15]
      enq_ptr_value <= 6'h0; // @[Counter.scala 98:11]
    end else if (do_enq) begin // @[Decoupled.scala 288:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 6'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 298:15]
      deq_ptr_value <= 6'h0; // @[Counter.scala 98:11]
    end else if (do_deq) begin // @[Decoupled.scala 292:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 278:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 278:27]
    end else if (io_flush) begin // @[Decoupled.scala 298:15]
      maybe_full <= 1'h0; // @[Decoupled.scala 301:16]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 295:27]
      maybe_full <= do_enq; // @[Decoupled.scala 296:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_io_deq_bits_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_io_deq_bits_MPORT_addr_pipe_0 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PISO(
  input        clock,
  input        reset,
  input        io_rd,
  input        io_wr,
  output       io_isEmpty,
  output       io_isAlmostEmpty,
  input  [7:0] io_din_0,
  input  [7:0] io_din_1,
  input  [7:0] io_din_2,
  input  [7:0] io_din_3,
  input  [7:0] io_din_4,
  input  [7:0] io_din_5,
  input  [7:0] io_din_6,
  input  [7:0] io_din_7,
  input  [7:0] io_din_8,
  input  [7:0] io_din_9,
  input  [7:0] io_din_10,
  input  [7:0] io_din_11,
  input  [7:0] io_din_12,
  input  [7:0] io_din_13,
  input  [7:0] io_din_14,
  input  [7:0] io_din_15,
  output [7:0] io_dout
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] pisoReg_0; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_1; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_2; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_3; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_4; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_5; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_6; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_7; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_8; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_9; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_10; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_11; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_12; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_13; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_14; // @[PISO.scala 61:20]
  reg [7:0] pisoReg_15; // @[PISO.scala 61:20]
  reg [4:0] pisoCounterReg; // @[PISO.scala 62:31]
  wire  pisoEmpty = pisoCounterReg == 5'h0; // @[PISO.scala 65:34]
  wire [4:0] _pisoCounterReg_T_1 = pisoCounterReg - 5'h1; // @[PISO.scala 74:38]
  assign io_isEmpty = pisoCounterReg == 5'h0; // @[PISO.scala 65:34]
  assign io_isAlmostEmpty = pisoCounterReg == 5'h1; // @[PISO.scala 66:40]
  assign io_dout = pisoReg_0; // @[PISO.scala 80:11]
  always @(posedge clock) begin
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_0 <= io_din_0; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_0 <= pisoReg_1; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_1 <= io_din_1; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_1 <= pisoReg_2; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_2 <= io_din_2; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_2 <= pisoReg_3; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_3 <= io_din_3; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_3 <= pisoReg_4; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_4 <= io_din_4; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_4 <= pisoReg_5; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_5 <= io_din_5; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_5 <= pisoReg_6; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_6 <= io_din_6; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_6 <= pisoReg_7; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_7 <= io_din_7; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_7 <= pisoReg_8; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_8 <= io_din_8; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_8 <= pisoReg_9; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_9 <= io_din_9; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_9 <= pisoReg_10; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_10 <= io_din_10; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_10 <= pisoReg_11; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_11 <= io_din_11; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_11 <= pisoReg_12; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_12 <= io_din_12; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_12 <= pisoReg_13; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_13 <= io_din_13; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_13 <= pisoReg_14; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_14 <= io_din_14; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_14 <= pisoReg_15; // @[PISO.scala 73:13]
    end
    if (io_wr) begin // @[PISO.scala 69:15]
      pisoReg_15 <= io_din_15; // @[PISO.scala 70:13]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoReg_15 <= pisoReg_0; // @[PISO.scala 73:13]
    end
    if (reset) begin // @[PISO.scala 62:31]
      pisoCounterReg <= 5'h0; // @[PISO.scala 62:31]
    end else if (io_wr) begin // @[PISO.scala 69:15]
      pisoCounterReg <= 5'h10; // @[PISO.scala 71:20]
    end else if (io_rd & ~pisoEmpty) begin // @[PISO.scala 72:35]
      pisoCounterReg <= _pisoCounterReg_T_1; // @[PISO.scala 74:20]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pisoReg_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  pisoReg_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  pisoReg_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  pisoReg_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  pisoReg_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  pisoReg_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  pisoReg_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  pisoReg_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  pisoReg_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  pisoReg_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  pisoReg_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  pisoReg_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  pisoReg_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  pisoReg_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  pisoReg_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  pisoReg_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  pisoCounterReg = _RAND_16[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SpriteBlitter(
  input         clock,
  input         reset,
  input         io_enable,
  output        io_busy,
  output        io_config_ready,
  input         io_config_valid,
  input  [1:0]  io_config_bits_sprite_priority,
  input  [5:0]  io_config_bits_sprite_colorCode,
  input         io_config_bits_sprite_hFlip,
  input         io_config_bits_sprite_vFlip,
  input  [17:0] io_config_bits_sprite_pos_x,
  input  [17:0] io_config_bits_sprite_pos_y,
  input  [7:0]  io_config_bits_sprite_cols,
  input  [7:0]  io_config_bits_sprite_rows,
  input  [15:0] io_config_bits_sprite_zoom_x,
  input  [15:0] io_config_bits_sprite_zoom_y,
  input         io_config_bits_hFlip,
  input  [8:0]  io_video_regs_size_x,
  input  [8:0]  io_video_regs_size_y,
  output        io_pixelData_ready,
  input         io_pixelData_valid,
  input  [7:0]  io_pixelData_bits_0,
  input  [7:0]  io_pixelData_bits_1,
  input  [7:0]  io_pixelData_bits_2,
  input  [7:0]  io_pixelData_bits_3,
  input  [7:0]  io_pixelData_bits_4,
  input  [7:0]  io_pixelData_bits_5,
  input  [7:0]  io_pixelData_bits_6,
  input  [7:0]  io_pixelData_bits_7,
  input  [7:0]  io_pixelData_bits_8,
  input  [7:0]  io_pixelData_bits_9,
  input  [7:0]  io_pixelData_bits_10,
  input  [7:0]  io_pixelData_bits_11,
  input  [7:0]  io_pixelData_bits_12,
  input  [7:0]  io_pixelData_bits_13,
  input  [7:0]  io_pixelData_bits_14,
  input  [7:0]  io_pixelData_bits_15,
  output        io_frameBuffer_wr,
  output [16:0] io_frameBuffer_addr,
  output [15:0] io_frameBuffer_din,
  input         io_frameBuffer_wait_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire  piso_clock; // @[SpriteBlitter.scala 74:20]
  wire  piso_reset; // @[SpriteBlitter.scala 74:20]
  wire  piso_io_rd; // @[SpriteBlitter.scala 74:20]
  wire  piso_io_wr; // @[SpriteBlitter.scala 74:20]
  wire  piso_io_isEmpty; // @[SpriteBlitter.scala 74:20]
  wire  piso_io_isAlmostEmpty; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_0; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_1; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_2; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_3; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_4; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_5; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_6; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_7; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_8; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_9; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_10; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_11; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_12; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_13; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_14; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_din_15; // @[SpriteBlitter.scala 74:20]
  wire [7:0] piso_io_dout; // @[SpriteBlitter.scala 74:20]
  reg  busyReg; // @[SpriteBlitter.scala 70:24]
  wire  _configReg_T = io_config_ready & io_config_valid; // @[Decoupled.scala 52:35]
  reg [1:0] configReg_sprite_priority; // @[Reg.scala 19:16]
  reg [5:0] configReg_sprite_colorCode; // @[Reg.scala 19:16]
  reg  configReg_sprite_hFlip; // @[Reg.scala 19:16]
  reg  configReg_sprite_vFlip; // @[Reg.scala 19:16]
  reg [17:0] configReg_sprite_pos_x; // @[Reg.scala 19:16]
  reg [17:0] configReg_sprite_pos_y; // @[Reg.scala 19:16]
  reg [7:0] configReg_sprite_cols; // @[Reg.scala 19:16]
  reg [7:0] configReg_sprite_rows; // @[Reg.scala 19:16]
  reg [15:0] configReg_sprite_zoom_x; // @[Reg.scala 19:16]
  reg [15:0] configReg_sprite_zoom_y; // @[Reg.scala 19:16]
  reg  configReg_hFlip; // @[Reg.scala 19:16]
  wire [11:0] vec_1_x = {configReg_sprite_cols, 4'h0}; // @[Vec2.scala 82:34]
  wire [11:0] vec_1_y = {configReg_sprite_rows, 4'h0}; // @[Vec2.scala 82:56]
  wire  _T_2 = ~piso_io_isEmpty; // @[SpriteBlitter.scala 84:81]
  wire  _T_4 = busyReg & ~piso_io_isEmpty & io_frameBuffer_wait_n; // @[SpriteBlitter.scala 84:92]
  reg [11:0] x; // @[Counter.scala 65:22]
  wire [11:0] _wrap_wrap_T_1 = vec_1_x - 12'h1; // @[Counter.scala 69:29]
  wire  wrap_wrap = x == _wrap_wrap_T_1 | vec_1_x == 12'h0; // @[Counter.scala 69:35]
  wire [11:0] _wrap_value_T_1 = x + 12'h1; // @[Counter.scala 70:20]
  wire  xWrap = _T_4 & wrap_wrap; // @[Counter.scala 93:{48,55}]
  reg [11:0] y; // @[Counter.scala 65:22]
  wire [11:0] _wrap_wrap_T_5 = vec_1_y - 12'h1; // @[Counter.scala 69:29]
  wire  wrap_wrap_1 = y == _wrap_wrap_T_5 | vec_1_y == 12'h0; // @[Counter.scala 69:35]
  wire [11:0] _wrap_value_T_3 = y + 12'h1; // @[Counter.scala 70:20]
  wire  yWrap = xWrap & wrap_wrap_1; // @[Counter.scala 93:{48,55}]
  wire [19:0] posReg_size_x = {vec_1_x, 8'h0}; // @[Vec2.scala 82:34]
  wire [19:0] posReg_size_y = {vec_1_y, 8'h0}; // @[Vec2.scala 82:56]
  wire [27:0] posReg_x = x * configReg_sprite_zoom_x; // @[SpriteBlitter.scala 140:19]
  wire [27:0] posReg_y = y * configReg_sprite_zoom_y; // @[SpriteBlitter.scala 141:19]
  wire [27:0] _GEN_31 = {{8'd0}, posReg_size_x}; // @[SpriteBlitter.scala 144:39]
  wire [27:0] _posReg_x__T_1 = _GEN_31 - posReg_x; // @[SpriteBlitter.scala 144:39]
  wire [27:0] _posReg_x__T_3 = _posReg_x__T_1 - 28'h100; // @[SpriteBlitter.scala 144:43]
  wire [27:0] _GEN_32 = {{8'd0}, posReg_size_y}; // @[SpriteBlitter.scala 145:39]
  wire [27:0] _posReg_y__T_1 = _GEN_32 - posReg_y; // @[SpriteBlitter.scala 145:39]
  wire [27:0] _posReg_y__T_3 = _posReg_y__T_1 - 28'h100; // @[SpriteBlitter.scala 145:43]
  wire [27:0] posReg_adjusted_vec_x = configReg_sprite_hFlip ? _posReg_x__T_3 : posReg_x; // @[Vec2.scala 159:16]
  wire [27:0] posReg_adjusted_vec_y = configReg_sprite_vFlip ? _posReg_y__T_3 : posReg_y; // @[Vec2.scala 160:16]
  wire [27:0] _GEN_33 = {{10{configReg_sprite_pos_x[17]}},configReg_sprite_pos_x}; // @[Vec2.scala 125:42]
  wire [27:0] posReg_adjusted_x = $signed(_GEN_33) + $signed(posReg_adjusted_vec_x); // @[Vec2.scala 125:42]
  wire [27:0] _GEN_34 = {{10{configReg_sprite_pos_y[17]}},configReg_sprite_pos_y}; // @[Vec2.scala 125:59]
  wire [27:0] posReg_adjusted_y = $signed(_GEN_34) + $signed(posReg_adjusted_vec_y); // @[Vec2.scala 125:59]
  wire [19:0] posReg_vec_1_x = posReg_adjusted_x[27:8]; // @[Vec2.scala 107:16]
  wire [19:0] posReg_vec_1_y = posReg_adjusted_y[27:8]; // @[Vec2.scala 108:16]
  reg [19:0] posReg__x; // @[Reg.scala 19:16]
  reg [19:0] posReg__y; // @[Reg.scala 19:16]
  reg [1:0] penReg_priority; // @[Reg.scala 19:16]
  reg [5:0] penReg_palette; // @[Reg.scala 19:16]
  reg [7:0] penReg_color; // @[Reg.scala 19:16]
  wire [7:0] pen_color = piso_io_dout; // @[PaletteEntry.scala 75:20 78:16]
  reg  validReg; // @[Reg.scala 19:16]
  wire [8:0] _visible_T_1 = io_video_regs_size_x - 9'h1; // @[SpriteBlitter.scala 184:37]
  wire [19:0] _GEN_35 = {{11'd0}, _visible_T_1}; // @[Util.scala 64:72]
  wire  _visible_T_3 = posReg__x <= _GEN_35; // @[Util.scala 64:72]
  wire [8:0] _visible_T_6 = io_video_regs_size_y - 9'h1; // @[SpriteBlitter.scala 184:79]
  wire [19:0] _GEN_36 = {{11'd0}, _visible_T_6}; // @[Util.scala 64:72]
  wire  _visible_T_8 = posReg__y <= _GEN_36; // @[Util.scala 64:72]
  wire  _visible_T_10 = _visible_T_3 & _visible_T_8; // @[SpriteBlitter.scala 184:44]
  wire  _visible_T_12 = penReg_color == 8'h0; // @[PaletteEntry.scala 63:35]
  wire  visible = _visible_T_10 & validReg & ~_visible_T_12; // @[SpriteBlitter.scala 96:76]
  wire  blitDone = xWrap & yWrap; // @[SpriteBlitter.scala 99:24]
  wire  _GEN_29 = blitDone ? 1'h0 : busyReg; // @[SpriteBlitter.scala 110:{65,75} 70:24]
  wire  _GEN_30 = _configReg_T | _GEN_29; // @[SpriteBlitter.scala 110:{24,34}]
  wire [19:0] _GEN_37 = {{11'd0}, io_video_regs_size_x}; // @[SpriteBlitter.scala 168:21]
  wire [19:0] _io_frameBuffer_addr_x__T_1 = _GEN_37 - posReg__x; // @[SpriteBlitter.scala 168:21]
  wire [19:0] io_frameBuffer_addr_x_ = _io_frameBuffer_addr_x__T_1 - 20'h1; // @[SpriteBlitter.scala 168:29]
  wire [19:0] _GEN_38 = {{11'd0}, io_video_regs_size_y}; // @[SpriteBlitter.scala 169:21]
  wire [19:0] _io_frameBuffer_addr_y__T_1 = _GEN_38 - posReg__y; // @[SpriteBlitter.scala 169:21]
  wire [19:0] io_frameBuffer_addr_y_ = _io_frameBuffer_addr_y__T_1 - 20'h1; // @[SpriteBlitter.scala 169:29]
  wire [28:0] _io_frameBuffer_addr_T = {io_frameBuffer_addr_y_, 9'h0}; // @[SpriteBlitter.scala 171:11]
  wire [28:0] _GEN_39 = {{9'd0}, io_frameBuffer_addr_x_}; // @[SpriteBlitter.scala 171:58]
  wire [28:0] _io_frameBuffer_addr_T_2 = _io_frameBuffer_addr_T + _GEN_39; // @[SpriteBlitter.scala 171:58]
  wire [28:0] _io_frameBuffer_addr_T_3 = {posReg__y, 9'h0}; // @[SpriteBlitter.scala 172:10]
  wire [28:0] _GEN_40 = {{9'd0}, posReg__x}; // @[SpriteBlitter.scala 172:57]
  wire [28:0] _io_frameBuffer_addr_T_5 = _io_frameBuffer_addr_T_3 + _GEN_40; // @[SpriteBlitter.scala 172:57]
  wire [28:0] _io_frameBuffer_addr_T_6 = configReg_hFlip ? _io_frameBuffer_addr_T_2 : _io_frameBuffer_addr_T_5; // @[SpriteBlitter.scala 170:8]
  wire [7:0] io_frameBuffer_din_hi = {penReg_priority,penReg_palette}; // @[SpriteBlitter.scala 118:32]
  PISO piso ( // @[SpriteBlitter.scala 74:20]
    .clock(piso_clock),
    .reset(piso_reset),
    .io_rd(piso_io_rd),
    .io_wr(piso_io_wr),
    .io_isEmpty(piso_io_isEmpty),
    .io_isAlmostEmpty(piso_io_isAlmostEmpty),
    .io_din_0(piso_io_din_0),
    .io_din_1(piso_io_din_1),
    .io_din_2(piso_io_din_2),
    .io_din_3(piso_io_din_3),
    .io_din_4(piso_io_din_4),
    .io_din_5(piso_io_din_5),
    .io_din_6(piso_io_din_6),
    .io_din_7(piso_io_din_7),
    .io_din_8(piso_io_din_8),
    .io_din_9(piso_io_din_9),
    .io_din_10(piso_io_din_10),
    .io_din_11(piso_io_din_11),
    .io_din_12(piso_io_din_12),
    .io_din_13(piso_io_din_13),
    .io_din_14(piso_io_din_14),
    .io_din_15(piso_io_din_15),
    .io_dout(piso_io_dout)
  );
  assign io_busy = busyReg; // @[SpriteBlitter.scala 119:11]
  assign io_config_ready = ~busyReg | blitDone; // @[SpriteBlitter.scala 103:30]
  assign io_pixelData_ready = io_frameBuffer_wait_n & (piso_io_isEmpty | piso_io_isAlmostEmpty); // @[SpriteBlitter.scala 107:46]
  assign io_frameBuffer_wr = io_enable & visible; // @[SpriteBlitter.scala 115:34]
  assign io_frameBuffer_addr = _io_frameBuffer_addr_T_6[16:0]; // @[SpriteBlitter.scala 116:23]
  assign io_frameBuffer_din = {io_frameBuffer_din_hi,penReg_color}; // @[SpriteBlitter.scala 118:32]
  assign piso_clock = clock;
  assign piso_reset = reset;
  assign piso_io_rd = busyReg & io_frameBuffer_wait_n; // @[SpriteBlitter.scala 75:25]
  assign piso_io_wr = io_pixelData_ready & io_pixelData_valid; // @[Decoupled.scala 52:35]
  assign piso_io_din_0 = io_pixelData_bits_0; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_1 = io_pixelData_bits_1; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_2 = io_pixelData_bits_2; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_3 = io_pixelData_bits_3; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_4 = io_pixelData_bits_4; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_5 = io_pixelData_bits_5; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_6 = io_pixelData_bits_6; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_7 = io_pixelData_bits_7; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_8 = io_pixelData_bits_8; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_9 = io_pixelData_bits_9; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_10 = io_pixelData_bits_10; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_11 = io_pixelData_bits_11; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_12 = io_pixelData_bits_12; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_13 = io_pixelData_bits_13; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_14 = io_pixelData_bits_14; // @[SpriteBlitter.scala 77:15]
  assign piso_io_din_15 = io_pixelData_bits_15; // @[SpriteBlitter.scala 77:15]
  always @(posedge clock) begin
    if (reset) begin // @[SpriteBlitter.scala 70:24]
      busyReg <= 1'h0; // @[SpriteBlitter.scala 70:24]
    end else begin
      busyReg <= _GEN_30;
    end
    if (_configReg_T) begin // @[Reg.scala 20:18]
      configReg_sprite_priority <= io_config_bits_sprite_priority; // @[Reg.scala 20:22]
    end
    if (_configReg_T) begin // @[Reg.scala 20:18]
      configReg_sprite_colorCode <= io_config_bits_sprite_colorCode; // @[Reg.scala 20:22]
    end
    if (_configReg_T) begin // @[Reg.scala 20:18]
      configReg_sprite_hFlip <= io_config_bits_sprite_hFlip; // @[Reg.scala 20:22]
    end
    if (_configReg_T) begin // @[Reg.scala 20:18]
      configReg_sprite_vFlip <= io_config_bits_sprite_vFlip; // @[Reg.scala 20:22]
    end
    if (_configReg_T) begin // @[Reg.scala 20:18]
      configReg_sprite_pos_x <= io_config_bits_sprite_pos_x; // @[Reg.scala 20:22]
    end
    if (_configReg_T) begin // @[Reg.scala 20:18]
      configReg_sprite_pos_y <= io_config_bits_sprite_pos_y; // @[Reg.scala 20:22]
    end
    if (_configReg_T) begin // @[Reg.scala 20:18]
      configReg_sprite_cols <= io_config_bits_sprite_cols; // @[Reg.scala 20:22]
    end
    if (_configReg_T) begin // @[Reg.scala 20:18]
      configReg_sprite_rows <= io_config_bits_sprite_rows; // @[Reg.scala 20:22]
    end
    if (_configReg_T) begin // @[Reg.scala 20:18]
      configReg_sprite_zoom_x <= io_config_bits_sprite_zoom_x; // @[Reg.scala 20:22]
    end
    if (_configReg_T) begin // @[Reg.scala 20:18]
      configReg_sprite_zoom_y <= io_config_bits_sprite_zoom_y; // @[Reg.scala 20:22]
    end
    if (_configReg_T) begin // @[Reg.scala 20:18]
      configReg_hFlip <= io_config_bits_hFlip; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[Counter.scala 65:22]
      x <= 12'h0; // @[Counter.scala 65:22]
    end else if (_T_4) begin // @[Counter.scala 93:48]
      if (wrap_wrap) begin // @[Counter.scala 71:16]
        x <= 12'h0; // @[Counter.scala 71:24]
      end else begin
        x <= _wrap_value_T_1; // @[Counter.scala 70:11]
      end
    end
    if (reset) begin // @[Counter.scala 65:22]
      y <= 12'h0; // @[Counter.scala 65:22]
    end else if (xWrap) begin // @[Counter.scala 93:48]
      if (wrap_wrap_1) begin // @[Counter.scala 71:16]
        y <= 12'h0; // @[Counter.scala 71:24]
      end else begin
        y <= _wrap_value_T_3; // @[Counter.scala 70:11]
      end
    end
    if (io_frameBuffer_wait_n) begin // @[Reg.scala 20:18]
      posReg__x <= posReg_vec_1_x; // @[Reg.scala 20:22]
    end
    if (io_frameBuffer_wait_n) begin // @[Reg.scala 20:18]
      posReg__y <= posReg_vec_1_y; // @[Reg.scala 20:22]
    end
    if (io_frameBuffer_wait_n) begin // @[Reg.scala 20:18]
      penReg_priority <= configReg_sprite_priority; // @[Reg.scala 20:22]
    end
    if (io_frameBuffer_wait_n) begin // @[Reg.scala 20:18]
      penReg_palette <= configReg_sprite_colorCode; // @[Reg.scala 20:22]
    end
    if (io_frameBuffer_wait_n) begin // @[Reg.scala 20:18]
      penReg_color <= pen_color; // @[Reg.scala 20:22]
    end
    if (io_frameBuffer_wait_n) begin // @[Reg.scala 20:18]
      validReg <= _T_2; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busyReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  configReg_sprite_priority = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  configReg_sprite_colorCode = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  configReg_sprite_hFlip = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  configReg_sprite_vFlip = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  configReg_sprite_pos_x = _RAND_5[17:0];
  _RAND_6 = {1{`RANDOM}};
  configReg_sprite_pos_y = _RAND_6[17:0];
  _RAND_7 = {1{`RANDOM}};
  configReg_sprite_cols = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  configReg_sprite_rows = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  configReg_sprite_zoom_x = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  configReg_sprite_zoom_y = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  configReg_hFlip = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  x = _RAND_12[11:0];
  _RAND_13 = {1{`RANDOM}};
  y = _RAND_13[11:0];
  _RAND_14 = {1{`RANDOM}};
  posReg__x = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  posReg__y = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  penReg_priority = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  penReg_palette = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  penReg_color = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  validReg = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SpriteDecoder(
  input         clock,
  input         reset,
  input  [1:0]  io_format,
  output        io_tileRom_ready,
  input         io_tileRom_valid,
  input  [63:0] io_tileRom_bits,
  input         io_pixelData_ready,
  output        io_pixelData_valid,
  output [7:0]  io_pixelData_bits_0,
  output [7:0]  io_pixelData_bits_1,
  output [7:0]  io_pixelData_bits_2,
  output [7:0]  io_pixelData_bits_3,
  output [7:0]  io_pixelData_bits_4,
  output [7:0]  io_pixelData_bits_5,
  output [7:0]  io_pixelData_bits_6,
  output [7:0]  io_pixelData_bits_7,
  output [7:0]  io_pixelData_bits_8,
  output [7:0]  io_pixelData_bits_9,
  output [7:0]  io_pixelData_bits_10,
  output [7:0]  io_pixelData_bits_11,
  output [7:0]  io_pixelData_bits_12,
  output [7:0]  io_pixelData_bits_13,
  output [7:0]  io_pixelData_bits_14,
  output [7:0]  io_pixelData_bits_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [127:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  is8BPP = io_format == 2'h3; // @[SpriteDecoder.scala 60:26]
  reg  pendingReg; // @[SpriteDecoder.scala 63:27]
  reg  validReg; // @[SpriteDecoder.scala 64:25]
  reg  toggleReg; // @[SpriteDecoder.scala 65:26]
  reg [127:0] dataReg; // @[SpriteDecoder.scala 66:20]
  wire  start = io_pixelData_ready & ~pendingReg; // @[SpriteDecoder.scala 69:34]
  wire  done = ~is8BPP | toggleReg; // @[SpriteDecoder.scala 70:22]
  wire [7:0] _bits_T_17 = {{4'd0}, dataReg[3:0]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_18 = {{4'd0}, dataReg[7:4]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_19 = {{4'd0}, dataReg[11:8]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_20 = {{4'd0}, dataReg[15:12]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_21 = {{4'd0}, dataReg[19:16]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_22 = {{4'd0}, dataReg[23:20]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_23 = {{4'd0}, dataReg[27:24]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_24 = {{4'd0}, dataReg[31:28]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_25 = {{4'd0}, dataReg[35:32]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_26 = {{4'd0}, dataReg[39:36]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_27 = {{4'd0}, dataReg[43:40]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_28 = {{4'd0}, dataReg[47:44]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_29 = {{4'd0}, dataReg[51:48]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_30 = {{4'd0}, dataReg[55:52]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_31 = {{4'd0}, dataReg[59:56]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_32 = {{4'd0}, dataReg[63:60]}; // @[SpriteDecoder.scala 113:17]
  wire [7:0] _bits_T_98 = {dataReg[67:64],dataReg[75:72]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_99 = {dataReg[71:68],dataReg[79:76]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_100 = {dataReg[83:80],dataReg[91:88]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_101 = {dataReg[87:84],dataReg[95:92]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_102 = {dataReg[99:96],dataReg[107:104]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_103 = {dataReg[103:100],dataReg[111:108]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_104 = {dataReg[115:112],dataReg[123:120]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_105 = {dataReg[119:116],dataReg[127:124]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_106 = {dataReg[3:0],dataReg[11:8]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_107 = {dataReg[7:4],dataReg[15:12]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_108 = {dataReg[19:16],dataReg[27:24]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_109 = {dataReg[23:20],dataReg[31:28]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_110 = {dataReg[35:32],dataReg[43:40]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_111 = {dataReg[39:36],dataReg[47:44]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_112 = {dataReg[51:48],dataReg[59:56]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_113 = {dataReg[55:52],dataReg[63:60]}; // @[Cat.scala 33:92]
  wire [7:0] _bits_T_115_0 = 2'h2 == io_format ? _bits_T_20 : _bits_T_17; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_1 = 2'h2 == io_format ? _bits_T_19 : _bits_T_18; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_2 = 2'h2 == io_format ? _bits_T_18 : _bits_T_19; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_3 = 2'h2 == io_format ? _bits_T_17 : _bits_T_20; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_4 = 2'h2 == io_format ? _bits_T_24 : _bits_T_21; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_5 = 2'h2 == io_format ? _bits_T_23 : _bits_T_22; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_6 = 2'h2 == io_format ? _bits_T_22 : _bits_T_23; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_7 = 2'h2 == io_format ? _bits_T_21 : _bits_T_24; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_8 = 2'h2 == io_format ? _bits_T_28 : _bits_T_25; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_9 = 2'h2 == io_format ? _bits_T_27 : _bits_T_26; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_10 = 2'h2 == io_format ? _bits_T_26 : _bits_T_27; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_11 = 2'h2 == io_format ? _bits_T_25 : _bits_T_28; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_12 = 2'h2 == io_format ? _bits_T_32 : _bits_T_29; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_13 = 2'h2 == io_format ? _bits_T_31 : _bits_T_30; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_14 = 2'h2 == io_format ? _bits_T_30 : _bits_T_31; // @[Mux.scala 81:58]
  wire [7:0] _bits_T_115_15 = 2'h2 == io_format ? _bits_T_29 : _bits_T_32; // @[Mux.scala 81:58]
  wire  _GEN_0 = start | pendingReg; // @[SpriteDecoder.scala 79:15 80:16 63:27]
  wire  _GEN_1 = start ? 1'h0 : validReg; // @[SpriteDecoder.scala 79:15 81:14 64:25]
  wire  _T = io_tileRom_ready & io_tileRom_valid; // @[Decoupled.scala 52:35]
  wire  _GEN_4 = done | _GEN_1; // @[SpriteDecoder.scala 87:16 89:16]
  wire [127:0] _dataReg_T_1 = {dataReg[63:0],io_tileRom_bits}; // @[SpriteDecoder.scala 91:57]
  assign io_tileRom_ready = pendingReg; // @[SpriteDecoder.scala 96:20]
  assign io_pixelData_valid = validReg; // @[SpriteDecoder.scala 97:22]
  assign io_pixelData_bits_0 = 2'h3 == io_format ? _bits_T_98 : _bits_T_115_0; // @[Mux.scala 81:58]
  assign io_pixelData_bits_1 = 2'h3 == io_format ? _bits_T_99 : _bits_T_115_1; // @[Mux.scala 81:58]
  assign io_pixelData_bits_2 = 2'h3 == io_format ? _bits_T_100 : _bits_T_115_2; // @[Mux.scala 81:58]
  assign io_pixelData_bits_3 = 2'h3 == io_format ? _bits_T_101 : _bits_T_115_3; // @[Mux.scala 81:58]
  assign io_pixelData_bits_4 = 2'h3 == io_format ? _bits_T_102 : _bits_T_115_4; // @[Mux.scala 81:58]
  assign io_pixelData_bits_5 = 2'h3 == io_format ? _bits_T_103 : _bits_T_115_5; // @[Mux.scala 81:58]
  assign io_pixelData_bits_6 = 2'h3 == io_format ? _bits_T_104 : _bits_T_115_6; // @[Mux.scala 81:58]
  assign io_pixelData_bits_7 = 2'h3 == io_format ? _bits_T_105 : _bits_T_115_7; // @[Mux.scala 81:58]
  assign io_pixelData_bits_8 = 2'h3 == io_format ? _bits_T_106 : _bits_T_115_8; // @[Mux.scala 81:58]
  assign io_pixelData_bits_9 = 2'h3 == io_format ? _bits_T_107 : _bits_T_115_9; // @[Mux.scala 81:58]
  assign io_pixelData_bits_10 = 2'h3 == io_format ? _bits_T_108 : _bits_T_115_10; // @[Mux.scala 81:58]
  assign io_pixelData_bits_11 = 2'h3 == io_format ? _bits_T_109 : _bits_T_115_11; // @[Mux.scala 81:58]
  assign io_pixelData_bits_12 = 2'h3 == io_format ? _bits_T_110 : _bits_T_115_12; // @[Mux.scala 81:58]
  assign io_pixelData_bits_13 = 2'h3 == io_format ? _bits_T_111 : _bits_T_115_13; // @[Mux.scala 81:58]
  assign io_pixelData_bits_14 = 2'h3 == io_format ? _bits_T_112 : _bits_T_115_14; // @[Mux.scala 81:58]
  assign io_pixelData_bits_15 = 2'h3 == io_format ? _bits_T_113 : _bits_T_115_15; // @[Mux.scala 81:58]
  always @(posedge clock) begin
    if (reset) begin // @[SpriteDecoder.scala 63:27]
      pendingReg <= 1'h0; // @[SpriteDecoder.scala 63:27]
    end else if (_T) begin // @[SpriteDecoder.scala 86:25]
      if (done) begin // @[SpriteDecoder.scala 87:16]
        pendingReg <= 1'h0; // @[SpriteDecoder.scala 88:18]
      end else begin
        pendingReg <= _GEN_0;
      end
    end else begin
      pendingReg <= _GEN_0;
    end
    if (reset) begin // @[SpriteDecoder.scala 64:25]
      validReg <= 1'h0; // @[SpriteDecoder.scala 64:25]
    end else if (_T) begin // @[SpriteDecoder.scala 86:25]
      validReg <= _GEN_4;
    end else if (start) begin // @[SpriteDecoder.scala 79:15]
      validReg <= 1'h0; // @[SpriteDecoder.scala 81:14]
    end
    if (reset) begin // @[SpriteDecoder.scala 65:26]
      toggleReg <= 1'h0; // @[SpriteDecoder.scala 65:26]
    end else if (_T) begin // @[SpriteDecoder.scala 86:25]
      toggleReg <= ~toggleReg; // @[SpriteDecoder.scala 92:15]
    end else if (start) begin // @[SpriteDecoder.scala 79:15]
      toggleReg <= 1'h0; // @[SpriteDecoder.scala 82:15]
    end
    if (_T) begin // @[SpriteDecoder.scala 86:25]
      dataReg <= _dataReg_T_1; // @[SpriteDecoder.scala 91:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pendingReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  validReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  toggleReg = _RAND_2[0:0];
  _RAND_3 = {4{`RANDOM}};
  dataReg = _RAND_3[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SpriteProcessor(
  input          clock,
  input          reset,
  input          io_ctrl_enable,
  input  [1:0]   io_ctrl_format,
  input          io_ctrl_start,
  input          io_ctrl_zoom,
  input  [1:0]   io_ctrl_regs_bank,
  input          io_ctrl_regs_fixed,
  input          io_ctrl_regs_hFlip,
  output         io_ctrl_vram_rd,
  output [11:0]  io_ctrl_vram_addr,
  input  [127:0] io_ctrl_vram_dout,
  output         io_ctrl_tileRom_rd,
  output [31:0]  io_ctrl_tileRom_addr,
  input  [63:0]  io_ctrl_tileRom_dout,
  input          io_ctrl_tileRom_wait_n,
  input          io_ctrl_tileRom_valid,
  output [7:0]   io_ctrl_tileRom_burstLength,
  input          io_ctrl_tileRom_burstDone,
  input  [8:0]   io_video_regs_size_x,
  input  [8:0]   io_video_regs_size_y,
  output         io_frameBuffer_wr,
  output [16:0]  io_frameBuffer_addr,
  output [15:0]  io_frameBuffer_din,
  input          io_frameBuffer_wait_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  fifo_clock; // @[SpriteProcessor.scala 92:20]
  wire  fifo_reset; // @[SpriteProcessor.scala 92:20]
  wire  fifo_io_enq_ready; // @[SpriteProcessor.scala 92:20]
  wire  fifo_io_enq_valid; // @[SpriteProcessor.scala 92:20]
  wire [63:0] fifo_io_enq_bits; // @[SpriteProcessor.scala 92:20]
  wire  fifo_io_deq_ready; // @[SpriteProcessor.scala 92:20]
  wire  fifo_io_deq_valid; // @[SpriteProcessor.scala 92:20]
  wire [63:0] fifo_io_deq_bits; // @[SpriteProcessor.scala 92:20]
  wire [6:0] fifo_io_count; // @[SpriteProcessor.scala 92:20]
  wire  fifo_io_flush; // @[SpriteProcessor.scala 92:20]
  wire  blitter_clock; // @[SpriteProcessor.scala 96:23]
  wire  blitter_reset; // @[SpriteProcessor.scala 96:23]
  wire  blitter_io_enable; // @[SpriteProcessor.scala 96:23]
  wire  blitter_io_busy; // @[SpriteProcessor.scala 96:23]
  wire  blitter_io_config_ready; // @[SpriteProcessor.scala 96:23]
  wire  blitter_io_config_valid; // @[SpriteProcessor.scala 96:23]
  wire [1:0] blitter_io_config_bits_sprite_priority; // @[SpriteProcessor.scala 96:23]
  wire [5:0] blitter_io_config_bits_sprite_colorCode; // @[SpriteProcessor.scala 96:23]
  wire  blitter_io_config_bits_sprite_hFlip; // @[SpriteProcessor.scala 96:23]
  wire  blitter_io_config_bits_sprite_vFlip; // @[SpriteProcessor.scala 96:23]
  wire [17:0] blitter_io_config_bits_sprite_pos_x; // @[SpriteProcessor.scala 96:23]
  wire [17:0] blitter_io_config_bits_sprite_pos_y; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_config_bits_sprite_cols; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_config_bits_sprite_rows; // @[SpriteProcessor.scala 96:23]
  wire [15:0] blitter_io_config_bits_sprite_zoom_x; // @[SpriteProcessor.scala 96:23]
  wire [15:0] blitter_io_config_bits_sprite_zoom_y; // @[SpriteProcessor.scala 96:23]
  wire  blitter_io_config_bits_hFlip; // @[SpriteProcessor.scala 96:23]
  wire [8:0] blitter_io_video_regs_size_x; // @[SpriteProcessor.scala 96:23]
  wire [8:0] blitter_io_video_regs_size_y; // @[SpriteProcessor.scala 96:23]
  wire  blitter_io_pixelData_ready; // @[SpriteProcessor.scala 96:23]
  wire  blitter_io_pixelData_valid; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_0; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_1; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_2; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_3; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_4; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_5; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_6; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_7; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_8; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_9; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_10; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_11; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_12; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_13; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_14; // @[SpriteProcessor.scala 96:23]
  wire [7:0] blitter_io_pixelData_bits_15; // @[SpriteProcessor.scala 96:23]
  wire  blitter_io_frameBuffer_wr; // @[SpriteProcessor.scala 96:23]
  wire [16:0] blitter_io_frameBuffer_addr; // @[SpriteProcessor.scala 96:23]
  wire [15:0] blitter_io_frameBuffer_din; // @[SpriteProcessor.scala 96:23]
  wire  blitter_io_frameBuffer_wait_n; // @[SpriteProcessor.scala 96:23]
  wire  decoder_clock; // @[SpriteProcessor.scala 101:23]
  wire  decoder_reset; // @[SpriteProcessor.scala 101:23]
  wire [1:0] decoder_io_format; // @[SpriteProcessor.scala 101:23]
  wire  decoder_io_tileRom_ready; // @[SpriteProcessor.scala 101:23]
  wire  decoder_io_tileRom_valid; // @[SpriteProcessor.scala 101:23]
  wire [63:0] decoder_io_tileRom_bits; // @[SpriteProcessor.scala 101:23]
  wire  decoder_io_pixelData_ready; // @[SpriteProcessor.scala 101:23]
  wire  decoder_io_pixelData_valid; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_0; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_1; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_2; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_3; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_4; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_5; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_6; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_7; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_8; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_9; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_10; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_11; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_12; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_13; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_14; // @[SpriteProcessor.scala 101:23]
  wire [7:0] decoder_io_pixelData_bits_15; // @[SpriteProcessor.scala 101:23]
  wire  is8BPP = io_ctrl_format == 2'h3; // @[SpriteProcessor.scala 73:31]
  wire [15:0] sprite_words_0 = io_ctrl_vram_dout[15:0]; // @[Util.scala 104:11]
  wire [15:0] sprite_words_1 = io_ctrl_vram_dout[31:16]; // @[Util.scala 104:11]
  wire [15:0] sprite_words_2 = io_ctrl_vram_dout[47:32]; // @[Util.scala 104:11]
  wire [15:0] sprite_words_3 = io_ctrl_vram_dout[63:48]; // @[Util.scala 104:11]
  wire [15:0] sprite_words_4 = io_ctrl_vram_dout[79:64]; // @[Util.scala 104:11]
  wire [15:0] sprite_words_5 = io_ctrl_vram_dout[95:80]; // @[Util.scala 104:11]
  wire [15:0] sprite_words_6 = io_ctrl_vram_dout[111:96]; // @[Util.scala 104:11]
  wire [1:0] sprite_sprite_priority = sprite_words_2[5:4]; // @[Sprite.scala 157:32]
  wire [5:0] sprite_sprite_colorCode = sprite_words_2[13:8]; // @[Sprite.scala 158:33]
  wire [17:0] sprite_sprite_code = {sprite_words_2[1:0],sprite_words_3}; // @[Sprite.scala 159:35]
  wire  sprite_sprite_hFlip = sprite_words_2[3]; // @[Sprite.scala 160:29]
  wire  sprite_sprite_vFlip = sprite_words_2[2]; // @[Sprite.scala 161:29]
  wire [17:0] sprite_sprite_pos_vec_x = {sprite_words_0,2'h0}; // @[Vec2.scala 159:16]
  wire [17:0] sprite_sprite_pos_vec_y = {sprite_words_1,2'h0}; // @[Vec2.scala 160:16]
  wire [17:0] sprite_sprite_pos_vec_1_x = {sprite_words_0[9:0],8'h0}; // @[Vec2.scala 159:16]
  wire [17:0] sprite_sprite_pos_vec_1_y = {sprite_words_1[9:0],8'h0}; // @[Vec2.scala 160:16]
  wire [7:0] sprite_sprite_cols = sprite_words_6[15:8]; // @[Sprite.scala 163:28]
  wire [7:0] sprite_sprite_rows = sprite_words_6[7:0]; // @[Sprite.scala 164:28]
  wire [1:0] sprite_sprite_1_priority = sprite_words_0[5:4]; // @[Sprite.scala 120:32]
  wire [5:0] sprite_sprite_1_colorCode = sprite_words_0[13:8]; // @[Sprite.scala 121:33]
  wire [17:0] sprite_sprite_1_code = {sprite_words_0[1:0],sprite_words_1}; // @[Sprite.scala 122:35]
  wire  sprite_sprite_1_hFlip = sprite_words_0[3]; // @[Sprite.scala 123:29]
  wire  sprite_sprite_1_vFlip = sprite_words_0[2]; // @[Sprite.scala 124:29]
  wire [17:0] sprite_sprite_pos_vec_2_x = {sprite_words_2,2'h0}; // @[Vec2.scala 159:16]
  wire [17:0] sprite_sprite_pos_vec_2_y = {sprite_words_3,2'h0}; // @[Vec2.scala 160:16]
  wire [17:0] sprite_sprite_pos_vec_3_x = {sprite_words_2[9:0],8'h0}; // @[Vec2.scala 159:16]
  wire [17:0] sprite_sprite_pos_vec_3_y = {sprite_words_3[9:0],8'h0}; // @[Vec2.scala 160:16]
  wire [7:0] sprite_sprite_1_cols = sprite_words_4[15:8]; // @[Sprite.scala 126:28]
  wire [7:0] sprite_sprite_1_rows = sprite_words_4[7:0]; // @[Sprite.scala 127:28]
  reg [2:0] stateReg; // @[SpriteProcessor.scala 82:25]
  wire  _spriteReg_T = stateReg == 3'h2; // @[SpriteProcessor.scala 83:46]
  reg [1:0] spriteReg_priority; // @[Reg.scala 19:16]
  reg [5:0] spriteReg_colorCode; // @[Reg.scala 19:16]
  reg [17:0] spriteReg_code; // @[Reg.scala 19:16]
  reg  spriteReg_hFlip; // @[Reg.scala 19:16]
  reg  spriteReg_vFlip; // @[Reg.scala 19:16]
  reg [17:0] spriteReg_pos_x; // @[Reg.scala 19:16]
  reg [17:0] spriteReg_pos_y; // @[Reg.scala 19:16]
  reg [7:0] spriteReg_cols; // @[Reg.scala 19:16]
  reg [7:0] spriteReg_rows; // @[Reg.scala 19:16]
  reg [15:0] spriteReg_zoom_x; // @[Reg.scala 19:16]
  reg [15:0] spriteReg_zoom_y; // @[Reg.scala 19:16]
  wire [15:0] _numTilesReg_T = spriteReg_cols * spriteReg_rows; // @[SpriteProcessor.scala 84:46]
  wire  _numTilesReg_T_1 = stateReg == 3'h3; // @[SpriteProcessor.scala 84:73]
  reg [15:0] numTilesReg; // @[Reg.scala 19:16]
  reg  readPendingReg; // @[SpriteProcessor.scala 85:31]
  wire  _T = stateReg == 3'h6; // @[SpriteProcessor.scala 88:80]
  reg [9:0] spriteCounter; // @[Counter.scala 40:34]
  wire  wrap_wrap = spriteCounter == 10'h3ff; // @[Counter.scala 45:24]
  wire [9:0] _wrap_value_T_1 = spriteCounter + 10'h1; // @[Counter.scala 46:22]
  wire  spriteCounterWrap = _T & wrap_wrap; // @[Counter.scala 86:{48,55}]
  reg [15:0] tileCounter; // @[Counter.scala 65:22]
  wire [15:0] _wrap_wrap_T_1 = numTilesReg - 16'h1; // @[Counter.scala 69:29]
  wire  wrap_wrap_1 = tileCounter == _wrap_wrap_T_1 | numTilesReg == 16'h0; // @[Counter.scala 69:35]
  wire [15:0] _wrap_value_T_3 = tileCounter + 16'h1; // @[Counter.scala 70:20]
  wire  _tileRomRead_T_1 = ~readPendingReg; // @[SpriteProcessor.scala 108:5]
  wire  _tileRomRead_T_2 = stateReg == 3'h5 & _tileRomRead_T_1; // @[SpriteProcessor.scala 107:48]
  wire  _tileRomRead_T_3 = fifo_io_count <= 7'h20; // @[SpriteProcessor.scala 109:19]
  wire  tileRomRead = _tileRomRead_T_2 & _tileRomRead_T_3; // @[SpriteProcessor.scala 108:21]
  wire  effectiveRead = tileRomRead & io_ctrl_tileRom_wait_n; // @[SpriteProcessor.scala 112:32]
  wire  tileCounterWrap = effectiveRead & wrap_wrap_1; // @[Counter.scala 93:{48,55}]
  wire [17:0] _GEN_51 = {{2'd0}, tileCounter}; // @[SpriteProcessor.scala 119:37]
  wire [17:0] _tileRomAddr_T_1 = spriteReg_code + _GEN_51; // @[SpriteProcessor.scala 119:37]
  wire [3:0] _tileRomAddr_T_2 = is8BPP ? 4'h8 : 4'h7; // @[SpriteProcessor.scala 119:58]
  wire [32:0] _GEN_0 = {{15'd0}, _tileRomAddr_T_1}; // @[SpriteProcessor.scala 119:52]
  wire [32:0] tileRomAddr = _GEN_0 << _tileRomAddr_T_2; // @[SpriteProcessor.scala 119:52]
  wire [5:0] tileRomBurstLength = is8BPP ? 6'h20 : 6'h10; // @[SpriteProcessor.scala 122:31]
  wire  _GEN_21 = effectiveRead | readPendingReg; // @[SpriteProcessor.scala 127:29 128:20 85:31]
  wire  _stateReg_T_2 = spriteReg_cols != 8'h0 & spriteReg_rows != 8'h0; // @[Sprite.scala 65:38]
  wire [2:0] _stateReg_T_3 = _stateReg_T_2 ? 3'h4 : 3'h6; // @[SpriteProcessor.scala 163:38]
  wire [2:0] _GEN_40 = blitter_io_config_ready ? 3'h5 : stateReg; // @[SpriteProcessor.scala 167:{37,48} 82:25]
  wire [2:0] _GEN_41 = tileCounterWrap ? 3'h6 : stateReg; // @[SpriteProcessor.scala 172:{29,40} 82:25]
  wire [2:0] _stateReg_T_4 = spriteCounterWrap ? 3'h7 : 3'h1; // @[SpriteProcessor.scala 177:22]
  wire [2:0] _GEN_42 = ~blitter_io_busy ? 3'h0 : stateReg; // @[SpriteProcessor.scala 182:{30,41} 82:25]
  wire [2:0] _GEN_43 = 3'h7 == stateReg ? _GEN_42 : stateReg; // @[SpriteProcessor.scala 150:20 82:25]
  wire [2:0] _GEN_44 = 3'h6 == stateReg ? _stateReg_T_4 : _GEN_43; // @[SpriteProcessor.scala 150:20 177:16]
  wire [2:0] _GEN_45 = 3'h5 == stateReg ? _GEN_41 : _GEN_44; // @[SpriteProcessor.scala 150:20]
  wire [2:0] _GEN_46 = 3'h4 == stateReg ? _GEN_40 : _GEN_45; // @[SpriteProcessor.scala 150:20]
  wire [2:0] _GEN_47 = 3'h3 == stateReg ? _stateReg_T_3 : _GEN_46; // @[SpriteProcessor.scala 150:20 163:32]
  Queue_1 fifo ( // @[SpriteProcessor.scala 92:20]
    .clock(fifo_clock),
    .reset(fifo_reset),
    .io_enq_ready(fifo_io_enq_ready),
    .io_enq_valid(fifo_io_enq_valid),
    .io_enq_bits(fifo_io_enq_bits),
    .io_deq_ready(fifo_io_deq_ready),
    .io_deq_valid(fifo_io_deq_valid),
    .io_deq_bits(fifo_io_deq_bits),
    .io_count(fifo_io_count),
    .io_flush(fifo_io_flush)
  );
  SpriteBlitter blitter ( // @[SpriteProcessor.scala 96:23]
    .clock(blitter_clock),
    .reset(blitter_reset),
    .io_enable(blitter_io_enable),
    .io_busy(blitter_io_busy),
    .io_config_ready(blitter_io_config_ready),
    .io_config_valid(blitter_io_config_valid),
    .io_config_bits_sprite_priority(blitter_io_config_bits_sprite_priority),
    .io_config_bits_sprite_colorCode(blitter_io_config_bits_sprite_colorCode),
    .io_config_bits_sprite_hFlip(blitter_io_config_bits_sprite_hFlip),
    .io_config_bits_sprite_vFlip(blitter_io_config_bits_sprite_vFlip),
    .io_config_bits_sprite_pos_x(blitter_io_config_bits_sprite_pos_x),
    .io_config_bits_sprite_pos_y(blitter_io_config_bits_sprite_pos_y),
    .io_config_bits_sprite_cols(blitter_io_config_bits_sprite_cols),
    .io_config_bits_sprite_rows(blitter_io_config_bits_sprite_rows),
    .io_config_bits_sprite_zoom_x(blitter_io_config_bits_sprite_zoom_x),
    .io_config_bits_sprite_zoom_y(blitter_io_config_bits_sprite_zoom_y),
    .io_config_bits_hFlip(blitter_io_config_bits_hFlip),
    .io_video_regs_size_x(blitter_io_video_regs_size_x),
    .io_video_regs_size_y(blitter_io_video_regs_size_y),
    .io_pixelData_ready(blitter_io_pixelData_ready),
    .io_pixelData_valid(blitter_io_pixelData_valid),
    .io_pixelData_bits_0(blitter_io_pixelData_bits_0),
    .io_pixelData_bits_1(blitter_io_pixelData_bits_1),
    .io_pixelData_bits_2(blitter_io_pixelData_bits_2),
    .io_pixelData_bits_3(blitter_io_pixelData_bits_3),
    .io_pixelData_bits_4(blitter_io_pixelData_bits_4),
    .io_pixelData_bits_5(blitter_io_pixelData_bits_5),
    .io_pixelData_bits_6(blitter_io_pixelData_bits_6),
    .io_pixelData_bits_7(blitter_io_pixelData_bits_7),
    .io_pixelData_bits_8(blitter_io_pixelData_bits_8),
    .io_pixelData_bits_9(blitter_io_pixelData_bits_9),
    .io_pixelData_bits_10(blitter_io_pixelData_bits_10),
    .io_pixelData_bits_11(blitter_io_pixelData_bits_11),
    .io_pixelData_bits_12(blitter_io_pixelData_bits_12),
    .io_pixelData_bits_13(blitter_io_pixelData_bits_13),
    .io_pixelData_bits_14(blitter_io_pixelData_bits_14),
    .io_pixelData_bits_15(blitter_io_pixelData_bits_15),
    .io_frameBuffer_wr(blitter_io_frameBuffer_wr),
    .io_frameBuffer_addr(blitter_io_frameBuffer_addr),
    .io_frameBuffer_din(blitter_io_frameBuffer_din),
    .io_frameBuffer_wait_n(blitter_io_frameBuffer_wait_n)
  );
  SpriteDecoder decoder ( // @[SpriteProcessor.scala 101:23]
    .clock(decoder_clock),
    .reset(decoder_reset),
    .io_format(decoder_io_format),
    .io_tileRom_ready(decoder_io_tileRom_ready),
    .io_tileRom_valid(decoder_io_tileRom_valid),
    .io_tileRom_bits(decoder_io_tileRom_bits),
    .io_pixelData_ready(decoder_io_pixelData_ready),
    .io_pixelData_valid(decoder_io_pixelData_valid),
    .io_pixelData_bits_0(decoder_io_pixelData_bits_0),
    .io_pixelData_bits_1(decoder_io_pixelData_bits_1),
    .io_pixelData_bits_2(decoder_io_pixelData_bits_2),
    .io_pixelData_bits_3(decoder_io_pixelData_bits_3),
    .io_pixelData_bits_4(decoder_io_pixelData_bits_4),
    .io_pixelData_bits_5(decoder_io_pixelData_bits_5),
    .io_pixelData_bits_6(decoder_io_pixelData_bits_6),
    .io_pixelData_bits_7(decoder_io_pixelData_bits_7),
    .io_pixelData_bits_8(decoder_io_pixelData_bits_8),
    .io_pixelData_bits_9(decoder_io_pixelData_bits_9),
    .io_pixelData_bits_10(decoder_io_pixelData_bits_10),
    .io_pixelData_bits_11(decoder_io_pixelData_bits_11),
    .io_pixelData_bits_12(decoder_io_pixelData_bits_12),
    .io_pixelData_bits_13(decoder_io_pixelData_bits_13),
    .io_pixelData_bits_14(decoder_io_pixelData_bits_14),
    .io_pixelData_bits_15(decoder_io_pixelData_bits_15)
  );
  assign io_ctrl_vram_rd = stateReg == 3'h1; // @[SpriteProcessor.scala 188:31]
  assign io_ctrl_vram_addr = {io_ctrl_regs_bank,spriteCounter}; // @[SpriteProcessor.scala 116:41]
  assign io_ctrl_tileRom_rd = _tileRomRead_T_2 & _tileRomRead_T_3; // @[SpriteProcessor.scala 108:21]
  assign io_ctrl_tileRom_addr = tileRomAddr[31:0]; // @[SpriteProcessor.scala 191:24]
  assign io_ctrl_tileRom_burstLength = {{2'd0}, tileRomBurstLength}; // @[SpriteProcessor.scala 192:31]
  assign io_frameBuffer_wr = blitter_io_frameBuffer_wr; // @[SpriteProcessor.scala 193:18]
  assign io_frameBuffer_addr = blitter_io_frameBuffer_addr; // @[SpriteProcessor.scala 193:18]
  assign io_frameBuffer_din = blitter_io_frameBuffer_din; // @[SpriteProcessor.scala 193:18]
  assign fifo_clock = clock;
  assign fifo_reset = reset;
  assign fifo_io_enq_valid = io_ctrl_tileRom_valid; // @[SpriteProcessor.scala 143:31 Decoupled.scala 65:20 74:20]
  assign fifo_io_enq_bits = io_ctrl_tileRom_dout; // @[SpriteProcessor.scala 143:31 Decoupled.scala 66:19]
  assign fifo_io_deq_ready = decoder_io_tileRom_ready; // @[SpriteProcessor.scala 103:22]
  assign fifo_io_flush = stateReg == 3'h0; // @[SpriteProcessor.scala 93:26]
  assign blitter_clock = clock;
  assign blitter_reset = reset;
  assign blitter_io_enable = io_ctrl_enable; // @[SpriteProcessor.scala 97:21]
  assign blitter_io_config_valid = stateReg == 3'h4; // @[SpriteProcessor.scala 132:17]
  assign blitter_io_config_bits_sprite_priority = spriteReg_priority; // @[SpriteProcessor.scala 133:22 134:19]
  assign blitter_io_config_bits_sprite_colorCode = spriteReg_colorCode; // @[SpriteProcessor.scala 133:22 134:19]
  assign blitter_io_config_bits_sprite_hFlip = spriteReg_hFlip; // @[SpriteProcessor.scala 133:22 134:19]
  assign blitter_io_config_bits_sprite_vFlip = spriteReg_vFlip; // @[SpriteProcessor.scala 133:22 134:19]
  assign blitter_io_config_bits_sprite_pos_x = spriteReg_pos_x; // @[SpriteProcessor.scala 133:22 134:19]
  assign blitter_io_config_bits_sprite_pos_y = spriteReg_pos_y; // @[SpriteProcessor.scala 133:22 134:19]
  assign blitter_io_config_bits_sprite_cols = spriteReg_cols; // @[SpriteProcessor.scala 133:22 134:19]
  assign blitter_io_config_bits_sprite_rows = spriteReg_rows; // @[SpriteProcessor.scala 133:22 134:19]
  assign blitter_io_config_bits_sprite_zoom_x = spriteReg_zoom_x; // @[SpriteProcessor.scala 133:22 134:19]
  assign blitter_io_config_bits_sprite_zoom_y = spriteReg_zoom_y; // @[SpriteProcessor.scala 133:22 134:19]
  assign blitter_io_config_bits_hFlip = io_ctrl_regs_hFlip; // @[SpriteProcessor.scala 133:22 135:18]
  assign blitter_io_video_regs_size_x = io_video_regs_size_x; // @[SpriteProcessor.scala 98:20]
  assign blitter_io_video_regs_size_y = io_video_regs_size_y; // @[SpriteProcessor.scala 98:20]
  assign blitter_io_pixelData_valid = decoder_io_pixelData_valid; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_0 = decoder_io_pixelData_bits_0; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_1 = decoder_io_pixelData_bits_1; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_2 = decoder_io_pixelData_bits_2; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_3 = decoder_io_pixelData_bits_3; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_4 = decoder_io_pixelData_bits_4; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_5 = decoder_io_pixelData_bits_5; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_6 = decoder_io_pixelData_bits_6; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_7 = decoder_io_pixelData_bits_7; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_8 = decoder_io_pixelData_bits_8; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_9 = decoder_io_pixelData_bits_9; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_10 = decoder_io_pixelData_bits_10; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_11 = decoder_io_pixelData_bits_11; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_12 = decoder_io_pixelData_bits_12; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_13 = decoder_io_pixelData_bits_13; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_14 = decoder_io_pixelData_bits_14; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_pixelData_bits_15 = decoder_io_pixelData_bits_15; // @[SpriteProcessor.scala 104:24]
  assign blitter_io_frameBuffer_wait_n = io_frameBuffer_wait_n; // @[SpriteProcessor.scala 193:18]
  assign decoder_clock = clock;
  assign decoder_reset = reset;
  assign decoder_io_format = io_ctrl_format; // @[SpriteProcessor.scala 102:21]
  assign decoder_io_tileRom_valid = fifo_io_deq_valid; // @[SpriteProcessor.scala 103:22]
  assign decoder_io_tileRom_bits = fifo_io_deq_bits; // @[SpriteProcessor.scala 103:22]
  assign decoder_io_pixelData_ready = blitter_io_pixelData_ready; // @[SpriteProcessor.scala 104:24]
  always @(posedge clock) begin
    if (reset) begin // @[SpriteProcessor.scala 82:25]
      stateReg <= 3'h0; // @[SpriteProcessor.scala 82:25]
    end else if (3'h0 == stateReg) begin // @[SpriteProcessor.scala 150:20]
      if (io_ctrl_start) begin // @[SpriteProcessor.scala 153:27]
        stateReg <= 3'h1; // @[SpriteProcessor.scala 153:38]
      end
    end else if (3'h1 == stateReg) begin // @[SpriteProcessor.scala 150:20]
      stateReg <= 3'h2; // @[SpriteProcessor.scala 157:31]
    end else if (3'h2 == stateReg) begin // @[SpriteProcessor.scala 150:20]
      stateReg <= 3'h3; // @[SpriteProcessor.scala 160:32]
    end else begin
      stateReg <= _GEN_47;
    end
    if (_spriteReg_T) begin // @[Reg.scala 20:18]
      if (io_ctrl_zoom) begin // @[Sprite.scala 94:8]
        spriteReg_priority <= sprite_sprite_priority;
      end else begin
        spriteReg_priority <= sprite_sprite_1_priority;
      end
    end
    if (_spriteReg_T) begin // @[Reg.scala 20:18]
      if (io_ctrl_zoom) begin // @[Sprite.scala 94:8]
        spriteReg_colorCode <= sprite_sprite_colorCode;
      end else begin
        spriteReg_colorCode <= sprite_sprite_1_colorCode;
      end
    end
    if (_spriteReg_T) begin // @[Reg.scala 20:18]
      if (io_ctrl_zoom) begin // @[Sprite.scala 94:8]
        spriteReg_code <= sprite_sprite_code;
      end else begin
        spriteReg_code <= sprite_sprite_1_code;
      end
    end
    if (_spriteReg_T) begin // @[Reg.scala 20:18]
      if (io_ctrl_zoom) begin // @[Sprite.scala 94:8]
        spriteReg_hFlip <= sprite_sprite_hFlip;
      end else begin
        spriteReg_hFlip <= sprite_sprite_1_hFlip;
      end
    end
    if (_spriteReg_T) begin // @[Reg.scala 20:18]
      if (io_ctrl_zoom) begin // @[Sprite.scala 94:8]
        spriteReg_vFlip <= sprite_sprite_vFlip;
      end else begin
        spriteReg_vFlip <= sprite_sprite_1_vFlip;
      end
    end
    if (_spriteReg_T) begin // @[Reg.scala 20:18]
      if (io_ctrl_zoom) begin // @[Sprite.scala 94:8]
        if (io_ctrl_regs_fixed) begin // @[Sprite.scala 178:73]
          spriteReg_pos_x <= sprite_sprite_pos_vec_x;
        end else begin
          spriteReg_pos_x <= sprite_sprite_pos_vec_1_x;
        end
      end else if (io_ctrl_regs_fixed) begin // @[Sprite.scala 178:73]
        spriteReg_pos_x <= sprite_sprite_pos_vec_2_x;
      end else begin
        spriteReg_pos_x <= sprite_sprite_pos_vec_3_x;
      end
    end
    if (_spriteReg_T) begin // @[Reg.scala 20:18]
      if (io_ctrl_zoom) begin // @[Sprite.scala 94:8]
        if (io_ctrl_regs_fixed) begin // @[Sprite.scala 178:73]
          spriteReg_pos_y <= sprite_sprite_pos_vec_y;
        end else begin
          spriteReg_pos_y <= sprite_sprite_pos_vec_1_y;
        end
      end else if (io_ctrl_regs_fixed) begin // @[Sprite.scala 178:73]
        spriteReg_pos_y <= sprite_sprite_pos_vec_2_y;
      end else begin
        spriteReg_pos_y <= sprite_sprite_pos_vec_3_y;
      end
    end
    if (_spriteReg_T) begin // @[Reg.scala 20:18]
      if (io_ctrl_zoom) begin // @[Sprite.scala 94:8]
        spriteReg_cols <= sprite_sprite_cols;
      end else begin
        spriteReg_cols <= sprite_sprite_1_cols;
      end
    end
    if (_spriteReg_T) begin // @[Reg.scala 20:18]
      if (io_ctrl_zoom) begin // @[Sprite.scala 94:8]
        spriteReg_rows <= sprite_sprite_rows;
      end else begin
        spriteReg_rows <= sprite_sprite_1_rows;
      end
    end
    if (_spriteReg_T) begin // @[Reg.scala 20:18]
      if (io_ctrl_zoom) begin // @[Sprite.scala 94:8]
        spriteReg_zoom_x <= sprite_words_4;
      end else begin
        spriteReg_zoom_x <= 16'h100;
      end
    end
    if (_spriteReg_T) begin // @[Reg.scala 20:18]
      if (io_ctrl_zoom) begin // @[Sprite.scala 94:8]
        spriteReg_zoom_y <= sprite_words_5;
      end else begin
        spriteReg_zoom_y <= 16'h100;
      end
    end
    if (_numTilesReg_T_1) begin // @[Reg.scala 20:18]
      numTilesReg <= _numTilesReg_T; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[SpriteProcessor.scala 85:31]
      readPendingReg <= 1'h0; // @[SpriteProcessor.scala 85:31]
    end else if (io_ctrl_tileRom_burstDone) begin // @[SpriteProcessor.scala 125:35]
      readPendingReg <= 1'h0; // @[SpriteProcessor.scala 126:20]
    end else begin
      readPendingReg <= _GEN_21;
    end
    if (reset) begin // @[Counter.scala 40:34]
      spriteCounter <= 10'h0; // @[Counter.scala 40:34]
    end else if (_T) begin // @[Counter.scala 86:48]
      spriteCounter <= _wrap_value_T_1; // @[Counter.scala 46:13]
    end
    if (reset) begin // @[Counter.scala 65:22]
      tileCounter <= 16'h0; // @[Counter.scala 65:22]
    end else if (effectiveRead) begin // @[Counter.scala 93:48]
      if (wrap_wrap_1) begin // @[Counter.scala 71:16]
        tileCounter <= 16'h0; // @[Counter.scala 71:24]
      end else begin
        tileCounter <= _wrap_value_T_3; // @[Counter.scala 70:11]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  spriteReg_priority = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  spriteReg_colorCode = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  spriteReg_code = _RAND_3[17:0];
  _RAND_4 = {1{`RANDOM}};
  spriteReg_hFlip = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  spriteReg_vFlip = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  spriteReg_pos_x = _RAND_6[17:0];
  _RAND_7 = {1{`RANDOM}};
  spriteReg_pos_y = _RAND_7[17:0];
  _RAND_8 = {1{`RANDOM}};
  spriteReg_cols = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  spriteReg_rows = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  spriteReg_zoom_x = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  spriteReg_zoom_y = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  numTilesReg = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  readPendingReg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  spriteCounter = _RAND_14[9:0];
  _RAND_15 = {1{`RANDOM}};
  tileCounter = _RAND_15[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LayerProcessor(
  input         clock,
  input         io_ctrl_enable,
  input  [1:0]  io_ctrl_format,
  input         io_ctrl_regs_tileSize,
  input         io_ctrl_regs_enable,
  input         io_ctrl_regs_flipX,
  input         io_ctrl_regs_flipY,
  input         io_ctrl_regs_rowScrollEnable,
  input         io_ctrl_regs_rowSelectEnable,
  input  [8:0]  io_ctrl_regs_scroll_x,
  input  [8:0]  io_ctrl_regs_scroll_y,
  output [11:0] io_ctrl_vram8x8_addr,
  input  [31:0] io_ctrl_vram8x8_dout,
  output [9:0]  io_ctrl_vram16x16_addr,
  input  [31:0] io_ctrl_vram16x16_dout,
  output [8:0]  io_ctrl_lineRam_addr,
  input  [31:0] io_ctrl_lineRam_dout,
  output        io_ctrl_tileRom_rd,
  output [31:0] io_ctrl_tileRom_addr,
  input  [63:0] io_ctrl_tileRom_dout,
  input         io_video_clockEnable,
  input  [8:0]  io_video_pos_x,
  input  [8:0]  io_video_pos_y,
  input         io_video_vBlank,
  input  [8:0]  io_video_regs_size_x,
  input  [8:0]  io_video_regs_size_y,
  input  [8:0]  io_spriteOffset_x,
  input  [8:0]  io_spriteOffset_y,
  output [1:0]  io_pen_priority,
  output [5:0]  io_pen_palette,
  output [7:0]  io_pen_color
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] lineEffectReg_words_0 = io_ctrl_lineRam_dout[15:0]; // @[Util.scala 104:11]
  wire [15:0] lineEffectReg_words_1 = io_ctrl_lineRam_dout[31:16]; // @[Util.scala 104:11]
  reg [8:0] lineEffectReg_rowSelect; // @[Reg.scala 19:16]
  reg [8:0] lineEffectReg_rowScroll; // @[Reg.scala 19:16]
  wire [8:0] lineEffectReg_lineEffect_rowSelect = lineEffectReg_words_1[8:0]; // @[LineEffect.scala 64:26 66:26]
  wire [8:0] lineEffectReg_lineEffect_rowScroll = lineEffectReg_words_0[8:0]; // @[LineEffect.scala 64:26 65:26]
  wire  layerEnable = io_ctrl_enable & io_ctrl_format != 2'h0 & io_ctrl_regs_enable; // @[LayerProcessor.scala 63:94]
  wire [4:0] layerOffset_x = io_ctrl_regs_tileSize ? 5'h12 : 5'ha; // @[LayerProcessor.scala 155:16]
  wire [4:0] _layerOffset_T_1 = layerOffset_x + 5'h1; // @[LayerProcessor.scala 158:30]
  wire [4:0] _layerOffset_T_2 = io_ctrl_regs_flipX ? _layerOffset_T_1 : layerOffset_x; // @[LayerProcessor.scala 158:10]
  wire [8:0] layerOffset__y = io_ctrl_regs_flipY ? 9'h1ef : 9'h1ee; // @[LayerProcessor.scala 159:10]
  wire [8:0] pos_normal_vec_x = io_video_pos_x + io_ctrl_regs_scroll_x; // @[Vec2.scala 73:42]
  wire [8:0] pos_normal_vec_y = io_video_pos_y + io_ctrl_regs_scroll_y; // @[Vec2.scala 73:59]
  wire [8:0] pos_normal_vec_1_x = pos_normal_vec_x - io_spriteOffset_x; // @[Vec2.scala 76:42]
  wire [8:0] pos_normal_vec_1_y = pos_normal_vec_y - io_spriteOffset_y; // @[Vec2.scala 76:59]
  wire [8:0] layerOffset__x = {{4'd0}, _layerOffset_T_2}; // @[Vec2.scala 106:19 107:11]
  wire [8:0] pos_normal_x = pos_normal_vec_1_x - layerOffset__x; // @[Vec2.scala 76:42]
  wire [8:0] pos_normal_y = pos_normal_vec_1_y - layerOffset__y; // @[Vec2.scala 76:59]
  wire [8:0] pos_flipped_vec_x = io_video_regs_size_x - io_video_pos_x; // @[Vec2.scala 76:42]
  wire [8:0] pos_flipped_vec_y = io_video_regs_size_y - io_video_pos_y; // @[Vec2.scala 76:59]
  wire [8:0] pos_flipped_vec_1_x = pos_flipped_vec_x + io_ctrl_regs_scroll_x; // @[Vec2.scala 73:42]
  wire [8:0] pos_flipped_vec_1_y = pos_flipped_vec_y + io_ctrl_regs_scroll_y; // @[Vec2.scala 73:59]
  wire [8:0] pos_flipped_vec_2_x = pos_flipped_vec_1_x - io_spriteOffset_x; // @[Vec2.scala 76:42]
  wire [8:0] pos_flipped_vec_2_y = pos_flipped_vec_1_y - io_spriteOffset_y; // @[Vec2.scala 76:59]
  wire [8:0] pos_flipped_x = pos_flipped_vec_2_x + layerOffset__x; // @[Vec2.scala 73:42]
  wire [8:0] pos_flipped_y = pos_flipped_vec_2_y + layerOffset__y; // @[Vec2.scala 73:59]
  wire [8:0] pos_x = io_ctrl_regs_flipX ? pos_flipped_x : pos_normal_x; // @[LayerProcessor.scala 78:10]
  wire [8:0] pos_y = io_ctrl_regs_flipY ? pos_flipped_y : pos_normal_y; // @[LayerProcessor.scala 79:10]
  wire [8:0] _pos__x_T = io_ctrl_regs_rowScrollEnable ? lineEffectReg_rowScroll : 9'h0; // @[LayerProcessor.scala 85:16]
  wire [8:0] pos__x = _pos__x_T + pos_x; // @[LayerProcessor.scala 85:77]
  wire [8:0] pos__y = io_ctrl_regs_rowSelectEnable ? lineEffectReg_rowSelect : pos_y; // @[LayerProcessor.scala 86:16]
  wire [3:0] tileOffset_x = io_ctrl_regs_tileSize ? pos__x[3:0] : {{1'd0}, pos__x[2:0]}; // @[LayerProcessor.scala 184:16]
  wire [3:0] tileOffset_y = io_ctrl_regs_tileSize ? pos__y[3:0] : {{1'd0}, pos__y[2:0]}; // @[LayerProcessor.scala 185:16]
  wire  _latchTile_T = tileOffset_x == 4'h5; // @[LayerProcessor.scala 95:18]
  wire  _latchTile_T_3 = io_ctrl_regs_tileSize ? tileOffset_x == 4'ha : tileOffset_x == 4'h2; // @[LayerProcessor.scala 96:8]
  wire  _latchTile_T_4 = io_ctrl_regs_flipX ? _latchTile_T : _latchTile_T_3; // @[LayerProcessor.scala 94:46]
  wire  latchTile = io_video_clockEnable & _latchTile_T_4; // @[LayerProcessor.scala 94:40]
  wire  _latchColor_T = tileOffset_x == 4'h0; // @[LayerProcessor.scala 99:18]
  wire  _latchColor_T_3 = io_ctrl_regs_tileSize ? tileOffset_x == 4'hf : tileOffset_x == 4'h7; // @[LayerProcessor.scala 100:8]
  wire  _latchColor_T_4 = io_ctrl_regs_flipX ? _latchColor_T : _latchColor_T_3; // @[LayerProcessor.scala 98:47]
  wire  latchColor = io_video_clockEnable & _latchColor_T_4; // @[LayerProcessor.scala 98:41]
  wire  _latchPix_T_1 = tileOffset_x[2:0] == 3'h0; // @[LayerProcessor.scala 103:24]
  wire  _latchPix_T_3 = tileOffset_x[2:0] == 3'h7; // @[LayerProcessor.scala 104:24]
  wire  _latchPix_T_4 = io_ctrl_regs_flipX ? _latchPix_T_1 : _latchPix_T_3; // @[LayerProcessor.scala 102:45]
  wire  latchPix = io_video_clockEnable & _latchPix_T_4; // @[LayerProcessor.scala 102:39]
  wire [8:0] _lineRamAddr_T_1 = pos_y + 9'h1; // @[LayerProcessor.scala 109:51]
  wire [8:0] _lineRamAddr_T_3 = pos_y - 9'h1; // @[LayerProcessor.scala 109:64]
  wire [4:0] _vramAddr_large_T_2 = io_ctrl_regs_flipX ? 5'h1f : 5'h1; // @[LayerProcessor.scala 171:50]
  wire [4:0] _vramAddr_large_T_4 = pos__x[8:4] + _vramAddr_large_T_2; // @[LayerProcessor.scala 171:45]
  wire [9:0] vramAddr_large = {pos__y[8:4],_vramAddr_large_T_4}; // @[LayerProcessor.scala 171:29]
  wire [5:0] _vramAddr_small_T_2 = io_ctrl_regs_flipX ? 6'h3f : 6'h1; // @[LayerProcessor.scala 172:50]
  wire [5:0] _vramAddr_small_T_4 = pos__x[8:3] + _vramAddr_small_T_2; // @[LayerProcessor.scala 172:45]
  wire [11:0] vramAddr_small = {pos__y[8:3],_vramAddr_small_T_4}; // @[LayerProcessor.scala 172:29]
  wire [11:0] vramAddr = io_ctrl_regs_tileSize ? {{2'd0}, vramAddr_large} : vramAddr_small; // @[LayerProcessor.scala 173:8]
  wire [15:0] tile_words_0 = io_ctrl_vram16x16_dout[15:0]; // @[Util.scala 104:11]
  wire [15:0] tile_words_1 = io_ctrl_vram16x16_dout[31:16]; // @[Util.scala 104:11]
  wire [1:0] tile_tile_priority = tile_words_0[15:14]; // @[Tile.scala 69:30]
  wire [5:0] tile_tile_colorCode = tile_words_0[13:8]; // @[Tile.scala 70:31]
  wire [15:0] tile_words_0_1 = io_ctrl_vram8x8_dout[15:0]; // @[Util.scala 104:11]
  wire [15:0] tile_words_1_1 = io_ctrl_vram8x8_dout[31:16]; // @[Util.scala 104:11]
  wire [1:0] tile_tile_1_priority = tile_words_0_1[15:14]; // @[Tile.scala 92:30]
  wire [5:0] tile_tile_1_colorCode = tile_words_0_1[13:8]; // @[Tile.scala 93:31]
  wire [17:0] tile_tile_1_code = {tile_words_0_1[1:0],tile_words_1_1}; // @[Tile.scala 94:33]
  wire [17:0] tile_tile_code = {{2'd0}, tile_words_1}; // @[Tile.scala 68:20 71:15]
  reg [1:0] tileReg_priority; // @[Reg.scala 19:16]
  reg [5:0] tileReg_colorCode; // @[Reg.scala 19:16]
  reg [17:0] tileReg_code; // @[Reg.scala 19:16]
  reg [1:0] priorityReg; // @[Reg.scala 19:16]
  reg [5:0] colorReg; // @[Reg.scala 19:16]
  wire  pixReg_word = tileOffset_y[0]; // @[LayerProcessor.scala 219:24]
  wire [31:0] pixReg_pixels_4BPP_bits = pixReg_word ? io_ctrl_tileRom_dout[31:0] : io_ctrl_tileRom_dout[63:32]; // @[LayerProcessor.scala 235:19]
  wire [7:0] pixReg_pixels_4BPP_0 = {{4'd0}, pixReg_pixels_4BPP_bits[31:28]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_1 = {{4'd0}, pixReg_pixels_4BPP_bits[27:24]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_2 = {{4'd0}, pixReg_pixels_4BPP_bits[23:20]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_3 = {{4'd0}, pixReg_pixels_4BPP_bits[19:16]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_4 = {{4'd0}, pixReg_pixels_4BPP_bits[15:12]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_5 = {{4'd0}, pixReg_pixels_4BPP_bits[11:8]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_6 = {{4'd0}, pixReg_pixels_4BPP_bits[7:4]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_7 = {{4'd0}, pixReg_pixels_4BPP_bits[3:0]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_8BPP_0 = {io_ctrl_tileRom_dout[55:52],io_ctrl_tileRom_dout[63:60]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_1 = {io_ctrl_tileRom_dout[51:48],io_ctrl_tileRom_dout[59:56]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_2 = {io_ctrl_tileRom_dout[39:36],io_ctrl_tileRom_dout[47:44]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_3 = {io_ctrl_tileRom_dout[35:32],io_ctrl_tileRom_dout[43:40]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_4 = {io_ctrl_tileRom_dout[23:20],io_ctrl_tileRom_dout[31:28]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_5 = {io_ctrl_tileRom_dout[19:16],io_ctrl_tileRom_dout[27:24]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_6 = {io_ctrl_tileRom_dout[7:4],io_ctrl_tileRom_dout[15:12]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_7 = {io_ctrl_tileRom_dout[3:0],io_ctrl_tileRom_dout[11:8]}; // @[Cat.scala 33:92]
  wire  _pixReg_T = io_ctrl_format == 2'h3; // @[LayerProcessor.scala 222:16]
  reg [7:0] pixReg_0; // @[Reg.scala 19:16]
  reg [7:0] pixReg_1; // @[Reg.scala 19:16]
  reg [7:0] pixReg_2; // @[Reg.scala 19:16]
  reg [7:0] pixReg_3; // @[Reg.scala 19:16]
  reg [7:0] pixReg_4; // @[Reg.scala 19:16]
  reg [7:0] pixReg_5; // @[Reg.scala 19:16]
  reg [7:0] pixReg_6; // @[Reg.scala 19:16]
  reg [7:0] pixReg_7; // @[Reg.scala 19:16]
  wire [7:0] _GEN_16 = 3'h1 == tileOffset_x[2:0] ? pixReg_1 : pixReg_0; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_17 = 3'h2 == tileOffset_x[2:0] ? pixReg_2 : _GEN_16; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_18 = 3'h3 == tileOffset_x[2:0] ? pixReg_3 : _GEN_17; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_19 = 3'h4 == tileOffset_x[2:0] ? pixReg_4 : _GEN_18; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_20 = 3'h5 == tileOffset_x[2:0] ? pixReg_5 : _GEN_19; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_21 = 3'h6 == tileOffset_x[2:0] ? pixReg_6 : _GEN_20; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] pen_color = 3'h7 == tileOffset_x[2:0] ? pixReg_7 : _GEN_21; // @[PaletteEntry.scala 78:{16,16}]
  wire  _io_ctrl_tileRom_addr_format8x8x4_T = ~io_ctrl_regs_tileSize; // @[LayerProcessor.scala 198:23]
  wire  _io_ctrl_tileRom_addr_format8x8x4_T_1 = io_ctrl_format == 2'h1; // @[LayerProcessor.scala 198:58]
  wire  io_ctrl_tileRom_addr_format8x8x4 = ~io_ctrl_regs_tileSize & io_ctrl_format == 2'h1; // @[LayerProcessor.scala 198:43]
  wire  io_ctrl_tileRom_addr_format8x8x8 = _io_ctrl_tileRom_addr_format8x8x4_T & _pixReg_T; // @[LayerProcessor.scala 199:43]
  wire  io_ctrl_tileRom_addr_format16x16x4 = io_ctrl_regs_tileSize & _io_ctrl_tileRom_addr_format8x8x4_T_1; // @[LayerProcessor.scala 200:44]
  wire  io_ctrl_tileRom_addr_format16x16x8 = io_ctrl_regs_tileSize & _pixReg_T; // @[LayerProcessor.scala 201:44]
  wire [22:0] _io_ctrl_tileRom_addr_T_2 = {tileReg_code,tileOffset_y[2:1],3'h0}; // @[LayerProcessor.scala 204:45]
  wire [23:0] _io_ctrl_tileRom_addr_T_5 = {tileReg_code,tileOffset_y[2:0],3'h0}; // @[LayerProcessor.scala 205:45]
  wire  _io_ctrl_tileRom_addr_T_9 = ~tileOffset_x[3]; // @[LayerProcessor.scala 206:47]
  wire [24:0] _io_ctrl_tileRom_addr_T_13 = {tileReg_code,tileOffset_y[3],_io_ctrl_tileRom_addr_T_9,tileOffset_y[2:1],3'h0
    }; // @[LayerProcessor.scala 206:78]
  wire [25:0] _io_ctrl_tileRom_addr_T_21 = {tileReg_code,tileOffset_y[3],_io_ctrl_tileRom_addr_T_9,tileOffset_y[2:0],3'h0
    }; // @[LayerProcessor.scala 207:78]
  wire [25:0] _io_ctrl_tileRom_addr_T_22 = io_ctrl_tileRom_addr_format16x16x8 ? _io_ctrl_tileRom_addr_T_21 : 26'h0; // @[Mux.scala 101:16]
  wire [25:0] _io_ctrl_tileRom_addr_T_23 = io_ctrl_tileRom_addr_format16x16x4 ? {{1'd0}, _io_ctrl_tileRom_addr_T_13} :
    _io_ctrl_tileRom_addr_T_22; // @[Mux.scala 101:16]
  wire [25:0] _io_ctrl_tileRom_addr_T_24 = io_ctrl_tileRom_addr_format8x8x8 ? {{2'd0}, _io_ctrl_tileRom_addr_T_5} :
    _io_ctrl_tileRom_addr_T_23; // @[Mux.scala 101:16]
  wire [25:0] _io_ctrl_tileRom_addr_T_25 = io_ctrl_tileRom_addr_format8x8x4 ? {{3'd0}, _io_ctrl_tileRom_addr_T_2} :
    _io_ctrl_tileRom_addr_T_24; // @[Mux.scala 101:16]
  assign io_ctrl_vram8x8_addr = io_ctrl_regs_tileSize ? {{2'd0}, vramAddr_large} : vramAddr_small; // @[LayerProcessor.scala 173:8]
  assign io_ctrl_vram16x16_addr = vramAddr[9:0]; // @[LayerProcessor.scala 135:26]
  assign io_ctrl_lineRam_addr = io_ctrl_regs_flipY ? _lineRamAddr_T_1 : _lineRamAddr_T_3; // @[LayerProcessor.scala 109:24]
  assign io_ctrl_tileRom_rd = layerEnable & ~io_video_vBlank; // @[LayerProcessor.scala 68:33]
  assign io_ctrl_tileRom_addr = {{6'd0}, _io_ctrl_tileRom_addr_T_25}; // @[LayerProcessor.scala 137:24]
  assign io_pen_priority = layerEnable ? priorityReg : 2'h0; // @[LayerProcessor.scala 138:16]
  assign io_pen_palette = layerEnable ? colorReg : 6'h0; // @[LayerProcessor.scala 138:16]
  assign io_pen_color = layerEnable ? pen_color : 8'h0; // @[LayerProcessor.scala 138:16]
  always @(posedge clock) begin
    if (io_video_clockEnable) begin // @[Reg.scala 20:18]
      lineEffectReg_rowSelect <= lineEffectReg_lineEffect_rowSelect; // @[Reg.scala 20:22]
    end
    if (io_video_clockEnable) begin // @[Reg.scala 20:18]
      lineEffectReg_rowScroll <= lineEffectReg_lineEffect_rowScroll; // @[Reg.scala 20:22]
    end
    if (latchTile) begin // @[Reg.scala 20:18]
      if (io_ctrl_regs_tileSize) begin // @[LayerProcessor.scala 115:17]
        tileReg_priority <= tile_tile_priority;
      end else begin
        tileReg_priority <= tile_tile_1_priority;
      end
    end
    if (latchTile) begin // @[Reg.scala 20:18]
      if (io_ctrl_regs_tileSize) begin // @[LayerProcessor.scala 115:17]
        tileReg_colorCode <= tile_tile_colorCode;
      end else begin
        tileReg_colorCode <= tile_tile_1_colorCode;
      end
    end
    if (latchTile) begin // @[Reg.scala 20:18]
      if (io_ctrl_regs_tileSize) begin // @[LayerProcessor.scala 115:17]
        tileReg_code <= tile_tile_code;
      end else begin
        tileReg_code <= tile_tile_1_code;
      end
    end
    if (latchColor) begin // @[Reg.scala 20:18]
      priorityReg <= tileReg_priority; // @[Reg.scala 20:22]
    end
    if (latchColor) begin // @[Reg.scala 20:18]
      colorReg <= tileReg_colorCode; // @[Reg.scala 20:22]
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_0 <= pixReg_pixels_8BPP_0;
      end else begin
        pixReg_0 <= pixReg_pixels_4BPP_0;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_1 <= pixReg_pixels_8BPP_1;
      end else begin
        pixReg_1 <= pixReg_pixels_4BPP_1;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_2 <= pixReg_pixels_8BPP_2;
      end else begin
        pixReg_2 <= pixReg_pixels_4BPP_2;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_3 <= pixReg_pixels_8BPP_3;
      end else begin
        pixReg_3 <= pixReg_pixels_4BPP_3;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_4 <= pixReg_pixels_8BPP_4;
      end else begin
        pixReg_4 <= pixReg_pixels_4BPP_4;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_5 <= pixReg_pixels_8BPP_5;
      end else begin
        pixReg_5 <= pixReg_pixels_4BPP_5;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_6 <= pixReg_pixels_8BPP_6;
      end else begin
        pixReg_6 <= pixReg_pixels_4BPP_6;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_7 <= pixReg_pixels_8BPP_7;
      end else begin
        pixReg_7 <= pixReg_pixels_4BPP_7;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lineEffectReg_rowSelect = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  lineEffectReg_rowScroll = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  tileReg_priority = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  tileReg_colorCode = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  tileReg_code = _RAND_4[17:0];
  _RAND_5 = {1{`RANDOM}};
  priorityReg = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  colorReg = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  pixReg_0 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  pixReg_1 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  pixReg_2 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  pixReg_3 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  pixReg_4 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  pixReg_5 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  pixReg_6 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  pixReg_7 = _RAND_14[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LayerProcessor_1(
  input         clock,
  input         io_ctrl_enable,
  input  [1:0]  io_ctrl_format,
  input         io_ctrl_regs_tileSize,
  input         io_ctrl_regs_enable,
  input         io_ctrl_regs_flipX,
  input         io_ctrl_regs_flipY,
  input         io_ctrl_regs_rowScrollEnable,
  input         io_ctrl_regs_rowSelectEnable,
  input  [8:0]  io_ctrl_regs_scroll_x,
  input  [8:0]  io_ctrl_regs_scroll_y,
  output [11:0] io_ctrl_vram8x8_addr,
  input  [31:0] io_ctrl_vram8x8_dout,
  output [9:0]  io_ctrl_vram16x16_addr,
  input  [31:0] io_ctrl_vram16x16_dout,
  output [8:0]  io_ctrl_lineRam_addr,
  input  [31:0] io_ctrl_lineRam_dout,
  output        io_ctrl_tileRom_rd,
  output [31:0] io_ctrl_tileRom_addr,
  input  [63:0] io_ctrl_tileRom_dout,
  input         io_video_clockEnable,
  input  [8:0]  io_video_pos_x,
  input  [8:0]  io_video_pos_y,
  input         io_video_vBlank,
  input  [8:0]  io_video_regs_size_x,
  input  [8:0]  io_video_regs_size_y,
  input  [8:0]  io_spriteOffset_x,
  input  [8:0]  io_spriteOffset_y,
  output [1:0]  io_pen_priority,
  output [5:0]  io_pen_palette,
  output [7:0]  io_pen_color
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] lineEffectReg_words_0 = io_ctrl_lineRam_dout[15:0]; // @[Util.scala 104:11]
  wire [15:0] lineEffectReg_words_1 = io_ctrl_lineRam_dout[31:16]; // @[Util.scala 104:11]
  reg [8:0] lineEffectReg_rowSelect; // @[Reg.scala 19:16]
  reg [8:0] lineEffectReg_rowScroll; // @[Reg.scala 19:16]
  wire [8:0] lineEffectReg_lineEffect_rowSelect = lineEffectReg_words_1[8:0]; // @[LineEffect.scala 64:26 66:26]
  wire [8:0] lineEffectReg_lineEffect_rowScroll = lineEffectReg_words_0[8:0]; // @[LineEffect.scala 64:26 65:26]
  wire  layerEnable = io_ctrl_enable & io_ctrl_format != 2'h0 & io_ctrl_regs_enable; // @[LayerProcessor.scala 63:94]
  wire [4:0] layerOffset_x = io_ctrl_regs_tileSize ? 5'h11 : 5'h9; // @[LayerProcessor.scala 155:16]
  wire [4:0] _layerOffset_T_1 = layerOffset_x + 5'h1; // @[LayerProcessor.scala 158:30]
  wire [4:0] _layerOffset_T_2 = io_ctrl_regs_flipX ? _layerOffset_T_1 : layerOffset_x; // @[LayerProcessor.scala 158:10]
  wire [8:0] layerOffset__y = io_ctrl_regs_flipY ? 9'h1ef : 9'h1ee; // @[LayerProcessor.scala 159:10]
  wire [8:0] pos_normal_vec_x = io_video_pos_x + io_ctrl_regs_scroll_x; // @[Vec2.scala 73:42]
  wire [8:0] pos_normal_vec_y = io_video_pos_y + io_ctrl_regs_scroll_y; // @[Vec2.scala 73:59]
  wire [8:0] pos_normal_vec_1_x = pos_normal_vec_x - io_spriteOffset_x; // @[Vec2.scala 76:42]
  wire [8:0] pos_normal_vec_1_y = pos_normal_vec_y - io_spriteOffset_y; // @[Vec2.scala 76:59]
  wire [8:0] layerOffset__x = {{4'd0}, _layerOffset_T_2}; // @[Vec2.scala 106:19 107:11]
  wire [8:0] pos_normal_x = pos_normal_vec_1_x - layerOffset__x; // @[Vec2.scala 76:42]
  wire [8:0] pos_normal_y = pos_normal_vec_1_y - layerOffset__y; // @[Vec2.scala 76:59]
  wire [8:0] pos_flipped_vec_x = io_video_regs_size_x - io_video_pos_x; // @[Vec2.scala 76:42]
  wire [8:0] pos_flipped_vec_y = io_video_regs_size_y - io_video_pos_y; // @[Vec2.scala 76:59]
  wire [8:0] pos_flipped_vec_1_x = pos_flipped_vec_x + io_ctrl_regs_scroll_x; // @[Vec2.scala 73:42]
  wire [8:0] pos_flipped_vec_1_y = pos_flipped_vec_y + io_ctrl_regs_scroll_y; // @[Vec2.scala 73:59]
  wire [8:0] pos_flipped_vec_2_x = pos_flipped_vec_1_x - io_spriteOffset_x; // @[Vec2.scala 76:42]
  wire [8:0] pos_flipped_vec_2_y = pos_flipped_vec_1_y - io_spriteOffset_y; // @[Vec2.scala 76:59]
  wire [8:0] pos_flipped_x = pos_flipped_vec_2_x + layerOffset__x; // @[Vec2.scala 73:42]
  wire [8:0] pos_flipped_y = pos_flipped_vec_2_y + layerOffset__y; // @[Vec2.scala 73:59]
  wire [8:0] pos_x = io_ctrl_regs_flipX ? pos_flipped_x : pos_normal_x; // @[LayerProcessor.scala 78:10]
  wire [8:0] pos_y = io_ctrl_regs_flipY ? pos_flipped_y : pos_normal_y; // @[LayerProcessor.scala 79:10]
  wire [8:0] _pos__x_T = io_ctrl_regs_rowScrollEnable ? lineEffectReg_rowScroll : 9'h0; // @[LayerProcessor.scala 85:16]
  wire [8:0] pos__x = _pos__x_T + pos_x; // @[LayerProcessor.scala 85:77]
  wire [8:0] pos__y = io_ctrl_regs_rowSelectEnable ? lineEffectReg_rowSelect : pos_y; // @[LayerProcessor.scala 86:16]
  wire [3:0] tileOffset_x = io_ctrl_regs_tileSize ? pos__x[3:0] : {{1'd0}, pos__x[2:0]}; // @[LayerProcessor.scala 184:16]
  wire [3:0] tileOffset_y = io_ctrl_regs_tileSize ? pos__y[3:0] : {{1'd0}, pos__y[2:0]}; // @[LayerProcessor.scala 185:16]
  wire  _latchTile_T = tileOffset_x == 4'h5; // @[LayerProcessor.scala 95:18]
  wire  _latchTile_T_3 = io_ctrl_regs_tileSize ? tileOffset_x == 4'ha : tileOffset_x == 4'h2; // @[LayerProcessor.scala 96:8]
  wire  _latchTile_T_4 = io_ctrl_regs_flipX ? _latchTile_T : _latchTile_T_3; // @[LayerProcessor.scala 94:46]
  wire  latchTile = io_video_clockEnable & _latchTile_T_4; // @[LayerProcessor.scala 94:40]
  wire  _latchColor_T = tileOffset_x == 4'h0; // @[LayerProcessor.scala 99:18]
  wire  _latchColor_T_3 = io_ctrl_regs_tileSize ? tileOffset_x == 4'hf : tileOffset_x == 4'h7; // @[LayerProcessor.scala 100:8]
  wire  _latchColor_T_4 = io_ctrl_regs_flipX ? _latchColor_T : _latchColor_T_3; // @[LayerProcessor.scala 98:47]
  wire  latchColor = io_video_clockEnable & _latchColor_T_4; // @[LayerProcessor.scala 98:41]
  wire  _latchPix_T_1 = tileOffset_x[2:0] == 3'h0; // @[LayerProcessor.scala 103:24]
  wire  _latchPix_T_3 = tileOffset_x[2:0] == 3'h7; // @[LayerProcessor.scala 104:24]
  wire  _latchPix_T_4 = io_ctrl_regs_flipX ? _latchPix_T_1 : _latchPix_T_3; // @[LayerProcessor.scala 102:45]
  wire  latchPix = io_video_clockEnable & _latchPix_T_4; // @[LayerProcessor.scala 102:39]
  wire [8:0] _lineRamAddr_T_1 = pos_y + 9'h1; // @[LayerProcessor.scala 109:51]
  wire [8:0] _lineRamAddr_T_3 = pos_y - 9'h1; // @[LayerProcessor.scala 109:64]
  wire [4:0] _vramAddr_large_T_2 = io_ctrl_regs_flipX ? 5'h1f : 5'h1; // @[LayerProcessor.scala 171:50]
  wire [4:0] _vramAddr_large_T_4 = pos__x[8:4] + _vramAddr_large_T_2; // @[LayerProcessor.scala 171:45]
  wire [9:0] vramAddr_large = {pos__y[8:4],_vramAddr_large_T_4}; // @[LayerProcessor.scala 171:29]
  wire [5:0] _vramAddr_small_T_2 = io_ctrl_regs_flipX ? 6'h3f : 6'h1; // @[LayerProcessor.scala 172:50]
  wire [5:0] _vramAddr_small_T_4 = pos__x[8:3] + _vramAddr_small_T_2; // @[LayerProcessor.scala 172:45]
  wire [11:0] vramAddr_small = {pos__y[8:3],_vramAddr_small_T_4}; // @[LayerProcessor.scala 172:29]
  wire [11:0] vramAddr = io_ctrl_regs_tileSize ? {{2'd0}, vramAddr_large} : vramAddr_small; // @[LayerProcessor.scala 173:8]
  wire [15:0] tile_words_0 = io_ctrl_vram16x16_dout[15:0]; // @[Util.scala 104:11]
  wire [15:0] tile_words_1 = io_ctrl_vram16x16_dout[31:16]; // @[Util.scala 104:11]
  wire [1:0] tile_tile_priority = tile_words_0[15:14]; // @[Tile.scala 69:30]
  wire [5:0] tile_tile_colorCode = tile_words_0[13:8]; // @[Tile.scala 70:31]
  wire [15:0] tile_words_0_1 = io_ctrl_vram8x8_dout[15:0]; // @[Util.scala 104:11]
  wire [15:0] tile_words_1_1 = io_ctrl_vram8x8_dout[31:16]; // @[Util.scala 104:11]
  wire [1:0] tile_tile_1_priority = tile_words_0_1[15:14]; // @[Tile.scala 92:30]
  wire [5:0] tile_tile_1_colorCode = tile_words_0_1[13:8]; // @[Tile.scala 93:31]
  wire [17:0] tile_tile_1_code = {tile_words_0_1[1:0],tile_words_1_1}; // @[Tile.scala 94:33]
  wire [17:0] tile_tile_code = {{2'd0}, tile_words_1}; // @[Tile.scala 68:20 71:15]
  reg [1:0] tileReg_priority; // @[Reg.scala 19:16]
  reg [5:0] tileReg_colorCode; // @[Reg.scala 19:16]
  reg [17:0] tileReg_code; // @[Reg.scala 19:16]
  reg [1:0] priorityReg; // @[Reg.scala 19:16]
  reg [5:0] colorReg; // @[Reg.scala 19:16]
  wire  pixReg_word = tileOffset_y[0]; // @[LayerProcessor.scala 219:24]
  wire [31:0] pixReg_pixels_4BPP_bits = pixReg_word ? io_ctrl_tileRom_dout[31:0] : io_ctrl_tileRom_dout[63:32]; // @[LayerProcessor.scala 235:19]
  wire [7:0] pixReg_pixels_4BPP_0 = {{4'd0}, pixReg_pixels_4BPP_bits[31:28]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_1 = {{4'd0}, pixReg_pixels_4BPP_bits[27:24]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_2 = {{4'd0}, pixReg_pixels_4BPP_bits[23:20]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_3 = {{4'd0}, pixReg_pixels_4BPP_bits[19:16]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_4 = {{4'd0}, pixReg_pixels_4BPP_bits[15:12]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_5 = {{4'd0}, pixReg_pixels_4BPP_bits[11:8]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_6 = {{4'd0}, pixReg_pixels_4BPP_bits[7:4]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_7 = {{4'd0}, pixReg_pixels_4BPP_bits[3:0]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_8BPP_0 = {io_ctrl_tileRom_dout[55:52],io_ctrl_tileRom_dout[63:60]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_1 = {io_ctrl_tileRom_dout[51:48],io_ctrl_tileRom_dout[59:56]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_2 = {io_ctrl_tileRom_dout[39:36],io_ctrl_tileRom_dout[47:44]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_3 = {io_ctrl_tileRom_dout[35:32],io_ctrl_tileRom_dout[43:40]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_4 = {io_ctrl_tileRom_dout[23:20],io_ctrl_tileRom_dout[31:28]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_5 = {io_ctrl_tileRom_dout[19:16],io_ctrl_tileRom_dout[27:24]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_6 = {io_ctrl_tileRom_dout[7:4],io_ctrl_tileRom_dout[15:12]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_7 = {io_ctrl_tileRom_dout[3:0],io_ctrl_tileRom_dout[11:8]}; // @[Cat.scala 33:92]
  wire  _pixReg_T = io_ctrl_format == 2'h3; // @[LayerProcessor.scala 222:16]
  reg [7:0] pixReg_0; // @[Reg.scala 19:16]
  reg [7:0] pixReg_1; // @[Reg.scala 19:16]
  reg [7:0] pixReg_2; // @[Reg.scala 19:16]
  reg [7:0] pixReg_3; // @[Reg.scala 19:16]
  reg [7:0] pixReg_4; // @[Reg.scala 19:16]
  reg [7:0] pixReg_5; // @[Reg.scala 19:16]
  reg [7:0] pixReg_6; // @[Reg.scala 19:16]
  reg [7:0] pixReg_7; // @[Reg.scala 19:16]
  wire [7:0] _GEN_16 = 3'h1 == tileOffset_x[2:0] ? pixReg_1 : pixReg_0; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_17 = 3'h2 == tileOffset_x[2:0] ? pixReg_2 : _GEN_16; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_18 = 3'h3 == tileOffset_x[2:0] ? pixReg_3 : _GEN_17; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_19 = 3'h4 == tileOffset_x[2:0] ? pixReg_4 : _GEN_18; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_20 = 3'h5 == tileOffset_x[2:0] ? pixReg_5 : _GEN_19; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_21 = 3'h6 == tileOffset_x[2:0] ? pixReg_6 : _GEN_20; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] pen_color = 3'h7 == tileOffset_x[2:0] ? pixReg_7 : _GEN_21; // @[PaletteEntry.scala 78:{16,16}]
  wire  _io_ctrl_tileRom_addr_format8x8x4_T = ~io_ctrl_regs_tileSize; // @[LayerProcessor.scala 198:23]
  wire  _io_ctrl_tileRom_addr_format8x8x4_T_1 = io_ctrl_format == 2'h1; // @[LayerProcessor.scala 198:58]
  wire  io_ctrl_tileRom_addr_format8x8x4 = ~io_ctrl_regs_tileSize & io_ctrl_format == 2'h1; // @[LayerProcessor.scala 198:43]
  wire  io_ctrl_tileRom_addr_format8x8x8 = _io_ctrl_tileRom_addr_format8x8x4_T & _pixReg_T; // @[LayerProcessor.scala 199:43]
  wire  io_ctrl_tileRom_addr_format16x16x4 = io_ctrl_regs_tileSize & _io_ctrl_tileRom_addr_format8x8x4_T_1; // @[LayerProcessor.scala 200:44]
  wire  io_ctrl_tileRom_addr_format16x16x8 = io_ctrl_regs_tileSize & _pixReg_T; // @[LayerProcessor.scala 201:44]
  wire [22:0] _io_ctrl_tileRom_addr_T_2 = {tileReg_code,tileOffset_y[2:1],3'h0}; // @[LayerProcessor.scala 204:45]
  wire [23:0] _io_ctrl_tileRom_addr_T_5 = {tileReg_code,tileOffset_y[2:0],3'h0}; // @[LayerProcessor.scala 205:45]
  wire  _io_ctrl_tileRom_addr_T_9 = ~tileOffset_x[3]; // @[LayerProcessor.scala 206:47]
  wire [24:0] _io_ctrl_tileRom_addr_T_13 = {tileReg_code,tileOffset_y[3],_io_ctrl_tileRom_addr_T_9,tileOffset_y[2:1],3'h0
    }; // @[LayerProcessor.scala 206:78]
  wire [25:0] _io_ctrl_tileRom_addr_T_21 = {tileReg_code,tileOffset_y[3],_io_ctrl_tileRom_addr_T_9,tileOffset_y[2:0],3'h0
    }; // @[LayerProcessor.scala 207:78]
  wire [25:0] _io_ctrl_tileRom_addr_T_22 = io_ctrl_tileRom_addr_format16x16x8 ? _io_ctrl_tileRom_addr_T_21 : 26'h0; // @[Mux.scala 101:16]
  wire [25:0] _io_ctrl_tileRom_addr_T_23 = io_ctrl_tileRom_addr_format16x16x4 ? {{1'd0}, _io_ctrl_tileRom_addr_T_13} :
    _io_ctrl_tileRom_addr_T_22; // @[Mux.scala 101:16]
  wire [25:0] _io_ctrl_tileRom_addr_T_24 = io_ctrl_tileRom_addr_format8x8x8 ? {{2'd0}, _io_ctrl_tileRom_addr_T_5} :
    _io_ctrl_tileRom_addr_T_23; // @[Mux.scala 101:16]
  wire [25:0] _io_ctrl_tileRom_addr_T_25 = io_ctrl_tileRom_addr_format8x8x4 ? {{3'd0}, _io_ctrl_tileRom_addr_T_2} :
    _io_ctrl_tileRom_addr_T_24; // @[Mux.scala 101:16]
  assign io_ctrl_vram8x8_addr = io_ctrl_regs_tileSize ? {{2'd0}, vramAddr_large} : vramAddr_small; // @[LayerProcessor.scala 173:8]
  assign io_ctrl_vram16x16_addr = vramAddr[9:0]; // @[LayerProcessor.scala 135:26]
  assign io_ctrl_lineRam_addr = io_ctrl_regs_flipY ? _lineRamAddr_T_1 : _lineRamAddr_T_3; // @[LayerProcessor.scala 109:24]
  assign io_ctrl_tileRom_rd = layerEnable & ~io_video_vBlank; // @[LayerProcessor.scala 68:33]
  assign io_ctrl_tileRom_addr = {{6'd0}, _io_ctrl_tileRom_addr_T_25}; // @[LayerProcessor.scala 137:24]
  assign io_pen_priority = layerEnable ? priorityReg : 2'h0; // @[LayerProcessor.scala 138:16]
  assign io_pen_palette = layerEnable ? colorReg : 6'h0; // @[LayerProcessor.scala 138:16]
  assign io_pen_color = layerEnable ? pen_color : 8'h0; // @[LayerProcessor.scala 138:16]
  always @(posedge clock) begin
    if (io_video_clockEnable) begin // @[Reg.scala 20:18]
      lineEffectReg_rowSelect <= lineEffectReg_lineEffect_rowSelect; // @[Reg.scala 20:22]
    end
    if (io_video_clockEnable) begin // @[Reg.scala 20:18]
      lineEffectReg_rowScroll <= lineEffectReg_lineEffect_rowScroll; // @[Reg.scala 20:22]
    end
    if (latchTile) begin // @[Reg.scala 20:18]
      if (io_ctrl_regs_tileSize) begin // @[LayerProcessor.scala 115:17]
        tileReg_priority <= tile_tile_priority;
      end else begin
        tileReg_priority <= tile_tile_1_priority;
      end
    end
    if (latchTile) begin // @[Reg.scala 20:18]
      if (io_ctrl_regs_tileSize) begin // @[LayerProcessor.scala 115:17]
        tileReg_colorCode <= tile_tile_colorCode;
      end else begin
        tileReg_colorCode <= tile_tile_1_colorCode;
      end
    end
    if (latchTile) begin // @[Reg.scala 20:18]
      if (io_ctrl_regs_tileSize) begin // @[LayerProcessor.scala 115:17]
        tileReg_code <= tile_tile_code;
      end else begin
        tileReg_code <= tile_tile_1_code;
      end
    end
    if (latchColor) begin // @[Reg.scala 20:18]
      priorityReg <= tileReg_priority; // @[Reg.scala 20:22]
    end
    if (latchColor) begin // @[Reg.scala 20:18]
      colorReg <= tileReg_colorCode; // @[Reg.scala 20:22]
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_0 <= pixReg_pixels_8BPP_0;
      end else begin
        pixReg_0 <= pixReg_pixels_4BPP_0;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_1 <= pixReg_pixels_8BPP_1;
      end else begin
        pixReg_1 <= pixReg_pixels_4BPP_1;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_2 <= pixReg_pixels_8BPP_2;
      end else begin
        pixReg_2 <= pixReg_pixels_4BPP_2;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_3 <= pixReg_pixels_8BPP_3;
      end else begin
        pixReg_3 <= pixReg_pixels_4BPP_3;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_4 <= pixReg_pixels_8BPP_4;
      end else begin
        pixReg_4 <= pixReg_pixels_4BPP_4;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_5 <= pixReg_pixels_8BPP_5;
      end else begin
        pixReg_5 <= pixReg_pixels_4BPP_5;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_6 <= pixReg_pixels_8BPP_6;
      end else begin
        pixReg_6 <= pixReg_pixels_4BPP_6;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_7 <= pixReg_pixels_8BPP_7;
      end else begin
        pixReg_7 <= pixReg_pixels_4BPP_7;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lineEffectReg_rowSelect = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  lineEffectReg_rowScroll = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  tileReg_priority = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  tileReg_colorCode = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  tileReg_code = _RAND_4[17:0];
  _RAND_5 = {1{`RANDOM}};
  priorityReg = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  colorReg = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  pixReg_0 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  pixReg_1 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  pixReg_2 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  pixReg_3 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  pixReg_4 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  pixReg_5 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  pixReg_6 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  pixReg_7 = _RAND_14[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LayerProcessor_2(
  input         clock,
  input         io_ctrl_enable,
  input  [1:0]  io_ctrl_format,
  input         io_ctrl_regs_tileSize,
  input         io_ctrl_regs_enable,
  input         io_ctrl_regs_flipX,
  input         io_ctrl_regs_flipY,
  input         io_ctrl_regs_rowScrollEnable,
  input         io_ctrl_regs_rowSelectEnable,
  input  [8:0]  io_ctrl_regs_scroll_x,
  input  [8:0]  io_ctrl_regs_scroll_y,
  output [11:0] io_ctrl_vram8x8_addr,
  input  [31:0] io_ctrl_vram8x8_dout,
  output [9:0]  io_ctrl_vram16x16_addr,
  input  [31:0] io_ctrl_vram16x16_dout,
  output [8:0]  io_ctrl_lineRam_addr,
  input  [31:0] io_ctrl_lineRam_dout,
  output        io_ctrl_tileRom_rd,
  output [31:0] io_ctrl_tileRom_addr,
  input  [63:0] io_ctrl_tileRom_dout,
  input         io_video_clockEnable,
  input  [8:0]  io_video_pos_x,
  input  [8:0]  io_video_pos_y,
  input         io_video_vBlank,
  input  [8:0]  io_video_regs_size_x,
  input  [8:0]  io_video_regs_size_y,
  input  [8:0]  io_spriteOffset_x,
  input  [8:0]  io_spriteOffset_y,
  output [1:0]  io_pen_priority,
  output [5:0]  io_pen_palette,
  output [7:0]  io_pen_color
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] lineEffectReg_words_0 = io_ctrl_lineRam_dout[15:0]; // @[Util.scala 104:11]
  wire [15:0] lineEffectReg_words_1 = io_ctrl_lineRam_dout[31:16]; // @[Util.scala 104:11]
  reg [8:0] lineEffectReg_rowSelect; // @[Reg.scala 19:16]
  reg [8:0] lineEffectReg_rowScroll; // @[Reg.scala 19:16]
  wire [8:0] lineEffectReg_lineEffect_rowSelect = lineEffectReg_words_1[8:0]; // @[LineEffect.scala 64:26 66:26]
  wire [8:0] lineEffectReg_lineEffect_rowScroll = lineEffectReg_words_0[8:0]; // @[LineEffect.scala 64:26 65:26]
  wire  layerEnable = io_ctrl_enable & io_ctrl_format != 2'h0 & io_ctrl_regs_enable; // @[LayerProcessor.scala 63:94]
  wire [4:0] layerOffset_x = io_ctrl_regs_tileSize ? 5'h10 : 5'h8; // @[LayerProcessor.scala 155:16]
  wire [4:0] _layerOffset_T_1 = layerOffset_x + 5'h1; // @[LayerProcessor.scala 158:30]
  wire [4:0] _layerOffset_T_2 = io_ctrl_regs_flipX ? _layerOffset_T_1 : layerOffset_x; // @[LayerProcessor.scala 158:10]
  wire [8:0] layerOffset__y = io_ctrl_regs_flipY ? 9'h1ef : 9'h1ee; // @[LayerProcessor.scala 159:10]
  wire [8:0] pos_normal_vec_x = io_video_pos_x + io_ctrl_regs_scroll_x; // @[Vec2.scala 73:42]
  wire [8:0] pos_normal_vec_y = io_video_pos_y + io_ctrl_regs_scroll_y; // @[Vec2.scala 73:59]
  wire [8:0] pos_normal_vec_1_x = pos_normal_vec_x - io_spriteOffset_x; // @[Vec2.scala 76:42]
  wire [8:0] pos_normal_vec_1_y = pos_normal_vec_y - io_spriteOffset_y; // @[Vec2.scala 76:59]
  wire [8:0] layerOffset__x = {{4'd0}, _layerOffset_T_2}; // @[Vec2.scala 106:19 107:11]
  wire [8:0] pos_normal_x = pos_normal_vec_1_x - layerOffset__x; // @[Vec2.scala 76:42]
  wire [8:0] pos_normal_y = pos_normal_vec_1_y - layerOffset__y; // @[Vec2.scala 76:59]
  wire [8:0] pos_flipped_vec_x = io_video_regs_size_x - io_video_pos_x; // @[Vec2.scala 76:42]
  wire [8:0] pos_flipped_vec_y = io_video_regs_size_y - io_video_pos_y; // @[Vec2.scala 76:59]
  wire [8:0] pos_flipped_vec_1_x = pos_flipped_vec_x + io_ctrl_regs_scroll_x; // @[Vec2.scala 73:42]
  wire [8:0] pos_flipped_vec_1_y = pos_flipped_vec_y + io_ctrl_regs_scroll_y; // @[Vec2.scala 73:59]
  wire [8:0] pos_flipped_vec_2_x = pos_flipped_vec_1_x - io_spriteOffset_x; // @[Vec2.scala 76:42]
  wire [8:0] pos_flipped_vec_2_y = pos_flipped_vec_1_y - io_spriteOffset_y; // @[Vec2.scala 76:59]
  wire [8:0] pos_flipped_x = pos_flipped_vec_2_x + layerOffset__x; // @[Vec2.scala 73:42]
  wire [8:0] pos_flipped_y = pos_flipped_vec_2_y + layerOffset__y; // @[Vec2.scala 73:59]
  wire [8:0] pos_x = io_ctrl_regs_flipX ? pos_flipped_x : pos_normal_x; // @[LayerProcessor.scala 78:10]
  wire [8:0] pos_y = io_ctrl_regs_flipY ? pos_flipped_y : pos_normal_y; // @[LayerProcessor.scala 79:10]
  wire [8:0] _pos__x_T = io_ctrl_regs_rowScrollEnable ? lineEffectReg_rowScroll : 9'h0; // @[LayerProcessor.scala 85:16]
  wire [8:0] pos__x = _pos__x_T + pos_x; // @[LayerProcessor.scala 85:77]
  wire [8:0] pos__y = io_ctrl_regs_rowSelectEnable ? lineEffectReg_rowSelect : pos_y; // @[LayerProcessor.scala 86:16]
  wire [3:0] tileOffset_x = io_ctrl_regs_tileSize ? pos__x[3:0] : {{1'd0}, pos__x[2:0]}; // @[LayerProcessor.scala 184:16]
  wire [3:0] tileOffset_y = io_ctrl_regs_tileSize ? pos__y[3:0] : {{1'd0}, pos__y[2:0]}; // @[LayerProcessor.scala 185:16]
  wire  _latchTile_T = tileOffset_x == 4'h5; // @[LayerProcessor.scala 95:18]
  wire  _latchTile_T_3 = io_ctrl_regs_tileSize ? tileOffset_x == 4'ha : tileOffset_x == 4'h2; // @[LayerProcessor.scala 96:8]
  wire  _latchTile_T_4 = io_ctrl_regs_flipX ? _latchTile_T : _latchTile_T_3; // @[LayerProcessor.scala 94:46]
  wire  latchTile = io_video_clockEnable & _latchTile_T_4; // @[LayerProcessor.scala 94:40]
  wire  _latchColor_T = tileOffset_x == 4'h0; // @[LayerProcessor.scala 99:18]
  wire  _latchColor_T_3 = io_ctrl_regs_tileSize ? tileOffset_x == 4'hf : tileOffset_x == 4'h7; // @[LayerProcessor.scala 100:8]
  wire  _latchColor_T_4 = io_ctrl_regs_flipX ? _latchColor_T : _latchColor_T_3; // @[LayerProcessor.scala 98:47]
  wire  latchColor = io_video_clockEnable & _latchColor_T_4; // @[LayerProcessor.scala 98:41]
  wire  _latchPix_T_1 = tileOffset_x[2:0] == 3'h0; // @[LayerProcessor.scala 103:24]
  wire  _latchPix_T_3 = tileOffset_x[2:0] == 3'h7; // @[LayerProcessor.scala 104:24]
  wire  _latchPix_T_4 = io_ctrl_regs_flipX ? _latchPix_T_1 : _latchPix_T_3; // @[LayerProcessor.scala 102:45]
  wire  latchPix = io_video_clockEnable & _latchPix_T_4; // @[LayerProcessor.scala 102:39]
  wire [8:0] _lineRamAddr_T_1 = pos_y + 9'h1; // @[LayerProcessor.scala 109:51]
  wire [8:0] _lineRamAddr_T_3 = pos_y - 9'h1; // @[LayerProcessor.scala 109:64]
  wire [4:0] _vramAddr_large_T_2 = io_ctrl_regs_flipX ? 5'h1f : 5'h1; // @[LayerProcessor.scala 171:50]
  wire [4:0] _vramAddr_large_T_4 = pos__x[8:4] + _vramAddr_large_T_2; // @[LayerProcessor.scala 171:45]
  wire [9:0] vramAddr_large = {pos__y[8:4],_vramAddr_large_T_4}; // @[LayerProcessor.scala 171:29]
  wire [5:0] _vramAddr_small_T_2 = io_ctrl_regs_flipX ? 6'h3f : 6'h1; // @[LayerProcessor.scala 172:50]
  wire [5:0] _vramAddr_small_T_4 = pos__x[8:3] + _vramAddr_small_T_2; // @[LayerProcessor.scala 172:45]
  wire [11:0] vramAddr_small = {pos__y[8:3],_vramAddr_small_T_4}; // @[LayerProcessor.scala 172:29]
  wire [11:0] vramAddr = io_ctrl_regs_tileSize ? {{2'd0}, vramAddr_large} : vramAddr_small; // @[LayerProcessor.scala 173:8]
  wire [15:0] tile_words_0 = io_ctrl_vram16x16_dout[15:0]; // @[Util.scala 104:11]
  wire [15:0] tile_words_1 = io_ctrl_vram16x16_dout[31:16]; // @[Util.scala 104:11]
  wire [1:0] tile_tile_priority = tile_words_0[15:14]; // @[Tile.scala 69:30]
  wire [5:0] tile_tile_colorCode = tile_words_0[13:8]; // @[Tile.scala 70:31]
  wire [15:0] tile_words_0_1 = io_ctrl_vram8x8_dout[15:0]; // @[Util.scala 104:11]
  wire [15:0] tile_words_1_1 = io_ctrl_vram8x8_dout[31:16]; // @[Util.scala 104:11]
  wire [1:0] tile_tile_1_priority = tile_words_0_1[15:14]; // @[Tile.scala 92:30]
  wire [5:0] tile_tile_1_colorCode = tile_words_0_1[13:8]; // @[Tile.scala 93:31]
  wire [17:0] tile_tile_1_code = {tile_words_0_1[1:0],tile_words_1_1}; // @[Tile.scala 94:33]
  wire [17:0] tile_tile_code = {{2'd0}, tile_words_1}; // @[Tile.scala 68:20 71:15]
  reg [1:0] tileReg_priority; // @[Reg.scala 19:16]
  reg [5:0] tileReg_colorCode; // @[Reg.scala 19:16]
  reg [17:0] tileReg_code; // @[Reg.scala 19:16]
  reg [1:0] priorityReg; // @[Reg.scala 19:16]
  reg [5:0] colorReg; // @[Reg.scala 19:16]
  wire  pixReg_word = tileOffset_y[0]; // @[LayerProcessor.scala 219:24]
  wire [31:0] pixReg_pixels_4BPP_bits = pixReg_word ? io_ctrl_tileRom_dout[31:0] : io_ctrl_tileRom_dout[63:32]; // @[LayerProcessor.scala 235:19]
  wire [7:0] pixReg_pixels_4BPP_0 = {{4'd0}, pixReg_pixels_4BPP_bits[31:28]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_1 = {{4'd0}, pixReg_pixels_4BPP_bits[27:24]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_2 = {{4'd0}, pixReg_pixels_4BPP_bits[23:20]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_3 = {{4'd0}, pixReg_pixels_4BPP_bits[19:16]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_4 = {{4'd0}, pixReg_pixels_4BPP_bits[15:12]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_5 = {{4'd0}, pixReg_pixels_4BPP_bits[11:8]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_6 = {{4'd0}, pixReg_pixels_4BPP_bits[7:4]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_4BPP_7 = {{4'd0}, pixReg_pixels_4BPP_bits[3:0]}; // @[LayerProcessor.scala 240:17]
  wire [7:0] pixReg_pixels_8BPP_0 = {io_ctrl_tileRom_dout[55:52],io_ctrl_tileRom_dout[63:60]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_1 = {io_ctrl_tileRom_dout[51:48],io_ctrl_tileRom_dout[59:56]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_2 = {io_ctrl_tileRom_dout[39:36],io_ctrl_tileRom_dout[47:44]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_3 = {io_ctrl_tileRom_dout[35:32],io_ctrl_tileRom_dout[43:40]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_4 = {io_ctrl_tileRom_dout[23:20],io_ctrl_tileRom_dout[31:28]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_5 = {io_ctrl_tileRom_dout[19:16],io_ctrl_tileRom_dout[27:24]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_6 = {io_ctrl_tileRom_dout[7:4],io_ctrl_tileRom_dout[15:12]}; // @[Cat.scala 33:92]
  wire [7:0] pixReg_pixels_8BPP_7 = {io_ctrl_tileRom_dout[3:0],io_ctrl_tileRom_dout[11:8]}; // @[Cat.scala 33:92]
  wire  _pixReg_T = io_ctrl_format == 2'h3; // @[LayerProcessor.scala 222:16]
  reg [7:0] pixReg_0; // @[Reg.scala 19:16]
  reg [7:0] pixReg_1; // @[Reg.scala 19:16]
  reg [7:0] pixReg_2; // @[Reg.scala 19:16]
  reg [7:0] pixReg_3; // @[Reg.scala 19:16]
  reg [7:0] pixReg_4; // @[Reg.scala 19:16]
  reg [7:0] pixReg_5; // @[Reg.scala 19:16]
  reg [7:0] pixReg_6; // @[Reg.scala 19:16]
  reg [7:0] pixReg_7; // @[Reg.scala 19:16]
  wire [7:0] _GEN_16 = 3'h1 == tileOffset_x[2:0] ? pixReg_1 : pixReg_0; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_17 = 3'h2 == tileOffset_x[2:0] ? pixReg_2 : _GEN_16; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_18 = 3'h3 == tileOffset_x[2:0] ? pixReg_3 : _GEN_17; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_19 = 3'h4 == tileOffset_x[2:0] ? pixReg_4 : _GEN_18; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_20 = 3'h5 == tileOffset_x[2:0] ? pixReg_5 : _GEN_19; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] _GEN_21 = 3'h6 == tileOffset_x[2:0] ? pixReg_6 : _GEN_20; // @[PaletteEntry.scala 78:{16,16}]
  wire [7:0] pen_color = 3'h7 == tileOffset_x[2:0] ? pixReg_7 : _GEN_21; // @[PaletteEntry.scala 78:{16,16}]
  wire  _io_ctrl_tileRom_addr_format8x8x4_T = ~io_ctrl_regs_tileSize; // @[LayerProcessor.scala 198:23]
  wire  _io_ctrl_tileRom_addr_format8x8x4_T_1 = io_ctrl_format == 2'h1; // @[LayerProcessor.scala 198:58]
  wire  io_ctrl_tileRom_addr_format8x8x4 = ~io_ctrl_regs_tileSize & io_ctrl_format == 2'h1; // @[LayerProcessor.scala 198:43]
  wire  io_ctrl_tileRom_addr_format8x8x8 = _io_ctrl_tileRom_addr_format8x8x4_T & _pixReg_T; // @[LayerProcessor.scala 199:43]
  wire  io_ctrl_tileRom_addr_format16x16x4 = io_ctrl_regs_tileSize & _io_ctrl_tileRom_addr_format8x8x4_T_1; // @[LayerProcessor.scala 200:44]
  wire  io_ctrl_tileRom_addr_format16x16x8 = io_ctrl_regs_tileSize & _pixReg_T; // @[LayerProcessor.scala 201:44]
  wire [22:0] _io_ctrl_tileRom_addr_T_2 = {tileReg_code,tileOffset_y[2:1],3'h0}; // @[LayerProcessor.scala 204:45]
  wire [23:0] _io_ctrl_tileRom_addr_T_5 = {tileReg_code,tileOffset_y[2:0],3'h0}; // @[LayerProcessor.scala 205:45]
  wire  _io_ctrl_tileRom_addr_T_9 = ~tileOffset_x[3]; // @[LayerProcessor.scala 206:47]
  wire [24:0] _io_ctrl_tileRom_addr_T_13 = {tileReg_code,tileOffset_y[3],_io_ctrl_tileRom_addr_T_9,tileOffset_y[2:1],3'h0
    }; // @[LayerProcessor.scala 206:78]
  wire [25:0] _io_ctrl_tileRom_addr_T_21 = {tileReg_code,tileOffset_y[3],_io_ctrl_tileRom_addr_T_9,tileOffset_y[2:0],3'h0
    }; // @[LayerProcessor.scala 207:78]
  wire [25:0] _io_ctrl_tileRom_addr_T_22 = io_ctrl_tileRom_addr_format16x16x8 ? _io_ctrl_tileRom_addr_T_21 : 26'h0; // @[Mux.scala 101:16]
  wire [25:0] _io_ctrl_tileRom_addr_T_23 = io_ctrl_tileRom_addr_format16x16x4 ? {{1'd0}, _io_ctrl_tileRom_addr_T_13} :
    _io_ctrl_tileRom_addr_T_22; // @[Mux.scala 101:16]
  wire [25:0] _io_ctrl_tileRom_addr_T_24 = io_ctrl_tileRom_addr_format8x8x8 ? {{2'd0}, _io_ctrl_tileRom_addr_T_5} :
    _io_ctrl_tileRom_addr_T_23; // @[Mux.scala 101:16]
  wire [25:0] _io_ctrl_tileRom_addr_T_25 = io_ctrl_tileRom_addr_format8x8x4 ? {{3'd0}, _io_ctrl_tileRom_addr_T_2} :
    _io_ctrl_tileRom_addr_T_24; // @[Mux.scala 101:16]
  assign io_ctrl_vram8x8_addr = io_ctrl_regs_tileSize ? {{2'd0}, vramAddr_large} : vramAddr_small; // @[LayerProcessor.scala 173:8]
  assign io_ctrl_vram16x16_addr = vramAddr[9:0]; // @[LayerProcessor.scala 135:26]
  assign io_ctrl_lineRam_addr = io_ctrl_regs_flipY ? _lineRamAddr_T_1 : _lineRamAddr_T_3; // @[LayerProcessor.scala 109:24]
  assign io_ctrl_tileRom_rd = layerEnable & ~io_video_vBlank; // @[LayerProcessor.scala 68:33]
  assign io_ctrl_tileRom_addr = {{6'd0}, _io_ctrl_tileRom_addr_T_25}; // @[LayerProcessor.scala 137:24]
  assign io_pen_priority = layerEnable ? priorityReg : 2'h0; // @[LayerProcessor.scala 138:16]
  assign io_pen_palette = layerEnable ? colorReg : 6'h0; // @[LayerProcessor.scala 138:16]
  assign io_pen_color = layerEnable ? pen_color : 8'h0; // @[LayerProcessor.scala 138:16]
  always @(posedge clock) begin
    if (io_video_clockEnable) begin // @[Reg.scala 20:18]
      lineEffectReg_rowSelect <= lineEffectReg_lineEffect_rowSelect; // @[Reg.scala 20:22]
    end
    if (io_video_clockEnable) begin // @[Reg.scala 20:18]
      lineEffectReg_rowScroll <= lineEffectReg_lineEffect_rowScroll; // @[Reg.scala 20:22]
    end
    if (latchTile) begin // @[Reg.scala 20:18]
      if (io_ctrl_regs_tileSize) begin // @[LayerProcessor.scala 115:17]
        tileReg_priority <= tile_tile_priority;
      end else begin
        tileReg_priority <= tile_tile_1_priority;
      end
    end
    if (latchTile) begin // @[Reg.scala 20:18]
      if (io_ctrl_regs_tileSize) begin // @[LayerProcessor.scala 115:17]
        tileReg_colorCode <= tile_tile_colorCode;
      end else begin
        tileReg_colorCode <= tile_tile_1_colorCode;
      end
    end
    if (latchTile) begin // @[Reg.scala 20:18]
      if (io_ctrl_regs_tileSize) begin // @[LayerProcessor.scala 115:17]
        tileReg_code <= tile_tile_code;
      end else begin
        tileReg_code <= tile_tile_1_code;
      end
    end
    if (latchColor) begin // @[Reg.scala 20:18]
      priorityReg <= tileReg_priority; // @[Reg.scala 20:22]
    end
    if (latchColor) begin // @[Reg.scala 20:18]
      colorReg <= tileReg_colorCode; // @[Reg.scala 20:22]
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_0 <= pixReg_pixels_8BPP_0;
      end else begin
        pixReg_0 <= pixReg_pixels_4BPP_0;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_1 <= pixReg_pixels_8BPP_1;
      end else begin
        pixReg_1 <= pixReg_pixels_4BPP_1;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_2 <= pixReg_pixels_8BPP_2;
      end else begin
        pixReg_2 <= pixReg_pixels_4BPP_2;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_3 <= pixReg_pixels_8BPP_3;
      end else begin
        pixReg_3 <= pixReg_pixels_4BPP_3;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_4 <= pixReg_pixels_8BPP_4;
      end else begin
        pixReg_4 <= pixReg_pixels_4BPP_4;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_5 <= pixReg_pixels_8BPP_5;
      end else begin
        pixReg_5 <= pixReg_pixels_4BPP_5;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_6 <= pixReg_pixels_8BPP_6;
      end else begin
        pixReg_6 <= pixReg_pixels_4BPP_6;
      end
    end
    if (latchPix) begin // @[Reg.scala 20:18]
      if (io_ctrl_format == 2'h3) begin // @[LayerProcessor.scala 222:8]
        pixReg_7 <= pixReg_pixels_8BPP_7;
      end else begin
        pixReg_7 <= pixReg_pixels_4BPP_7;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lineEffectReg_rowSelect = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  lineEffectReg_rowScroll = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  tileReg_priority = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  tileReg_colorCode = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  tileReg_code = _RAND_4[17:0];
  _RAND_5 = {1{`RANDOM}};
  priorityReg = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  colorReg = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  pixReg_0 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  pixReg_1 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  pixReg_2 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  pixReg_3 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  pixReg_4 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  pixReg_5 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  pixReg_6 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  pixReg_7 = _RAND_14[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ColorMixer(
  input         clock,
  input  [8:0]  io_gameConfig_granularity,
  input  [1:0]  io_gameConfig_layer_0_paletteBank,
  input  [1:0]  io_gameConfig_layer_1_paletteBank,
  input  [1:0]  io_gameConfig_layer_2_paletteBank,
  input  [1:0]  io_spritePen_priority,
  input  [5:0]  io_spritePen_palette,
  input  [7:0]  io_spritePen_color,
  input  [1:0]  io_layer0Pen_priority,
  input  [5:0]  io_layer0Pen_palette,
  input  [7:0]  io_layer0Pen_color,
  input  [1:0]  io_layer1Pen_priority,
  input  [5:0]  io_layer1Pen_palette,
  input  [7:0]  io_layer1Pen_color,
  input  [1:0]  io_layer2Pen_priority,
  input  [5:0]  io_layer2Pen_palette,
  input  [7:0]  io_layer2Pen_color,
  output [14:0] io_paletteRam_addr,
  input  [15:0] io_paletteRam_dout,
  output [15:0] io_dout
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _index_T = io_spritePen_color != 8'h0; // @[ColorMixer.scala 116:24]
  wire  _index_T_2 = io_spritePen_color != 8'h0 & io_spritePen_priority == 2'h0; // @[ColorMixer.scala 116:32]
  wire  _index_T_5 = _index_T & io_spritePen_priority == 2'h1; // @[ColorMixer.scala 117:32]
  wire  _index_T_8 = _index_T & io_spritePen_priority == 2'h2; // @[ColorMixer.scala 118:32]
  wire  _index_T_11 = _index_T & io_spritePen_priority == 2'h3; // @[ColorMixer.scala 119:32]
  wire  _index_T_12 = io_layer0Pen_color != 8'h0; // @[ColorMixer.scala 123:24]
  wire  _index_T_14 = io_layer0Pen_color != 8'h0 & io_layer0Pen_priority == 2'h0; // @[ColorMixer.scala 123:32]
  wire  _index_T_17 = _index_T_12 & io_layer0Pen_priority == 2'h1; // @[ColorMixer.scala 124:32]
  wire  _index_T_20 = _index_T_12 & io_layer0Pen_priority == 2'h2; // @[ColorMixer.scala 125:32]
  wire  _index_T_23 = _index_T_12 & io_layer0Pen_priority == 2'h3; // @[ColorMixer.scala 126:32]
  wire  _index_T_24 = io_layer1Pen_color != 8'h0; // @[ColorMixer.scala 130:24]
  wire  _index_T_26 = io_layer1Pen_color != 8'h0 & io_layer1Pen_priority == 2'h0; // @[ColorMixer.scala 130:32]
  wire  _index_T_29 = _index_T_24 & io_layer1Pen_priority == 2'h1; // @[ColorMixer.scala 131:32]
  wire  _index_T_32 = _index_T_24 & io_layer1Pen_priority == 2'h2; // @[ColorMixer.scala 132:32]
  wire  _index_T_35 = _index_T_24 & io_layer1Pen_priority == 2'h3; // @[ColorMixer.scala 133:32]
  wire  _index_T_36 = io_layer2Pen_color != 8'h0; // @[ColorMixer.scala 137:24]
  wire  _index_T_38 = io_layer2Pen_color != 8'h0 & io_layer2Pen_priority == 2'h0; // @[ColorMixer.scala 137:32]
  wire  _index_T_41 = _index_T_36 & io_layer2Pen_priority == 2'h1; // @[ColorMixer.scala 138:32]
  wire  _index_T_44 = _index_T_36 & io_layer2Pen_priority == 2'h2; // @[ColorMixer.scala 139:32]
  wire  _index_T_47 = _index_T_36 & io_layer2Pen_priority == 2'h3; // @[ColorMixer.scala 140:32]
  wire [1:0] _index_T_49 = _index_T_14 ? 2'h2 : {{1'd0}, _index_T_2}; // @[Mux.scala 101:16]
  wire [2:0] _index_T_50 = _index_T_26 ? 3'h4 : {{1'd0}, _index_T_49}; // @[Mux.scala 101:16]
  wire [3:0] _index_T_51 = _index_T_38 ? 4'h8 : {{1'd0}, _index_T_50}; // @[Mux.scala 101:16]
  wire [3:0] _index_T_52 = _index_T_5 ? 4'h1 : _index_T_51; // @[Mux.scala 101:16]
  wire [3:0] _index_T_53 = _index_T_17 ? 4'h2 : _index_T_52; // @[Mux.scala 101:16]
  wire [3:0] _index_T_54 = _index_T_29 ? 4'h4 : _index_T_53; // @[Mux.scala 101:16]
  wire [3:0] _index_T_55 = _index_T_41 ? 4'h8 : _index_T_54; // @[Mux.scala 101:16]
  wire [3:0] _index_T_56 = _index_T_8 ? 4'h1 : _index_T_55; // @[Mux.scala 101:16]
  wire [3:0] _index_T_57 = _index_T_20 ? 4'h2 : _index_T_56; // @[Mux.scala 101:16]
  wire [3:0] _index_T_58 = _index_T_32 ? 4'h4 : _index_T_57; // @[Mux.scala 101:16]
  wire [3:0] _index_T_59 = _index_T_44 ? 4'h8 : _index_T_58; // @[Mux.scala 101:16]
  wire [3:0] _index_T_60 = _index_T_11 ? 4'h1 : _index_T_59; // @[Mux.scala 101:16]
  wire [3:0] _index_T_61 = _index_T_23 ? 4'h2 : _index_T_60; // @[Mux.scala 101:16]
  wire [3:0] _index_T_62 = _index_T_35 ? 4'h4 : _index_T_61; // @[Mux.scala 101:16]
  wire [3:0] index = _index_T_47 ? 4'h8 : _index_T_62; // @[Mux.scala 101:16]
  wire [14:0] _paletteRamAddr_T_9 = 9'h10 == io_gameConfig_granularity ? 15'h3f0 : 15'h3f00; // @[Mux.scala 81:58]
  wire [14:0] _paletteRamAddr_T_11 = 9'h40 == io_gameConfig_granularity ? 15'hfc0 : _paletteRamAddr_T_9; // @[Mux.scala 81:58]
  wire [14:0] _paletteRamAddr_T_13 = {1'h0,io_spritePen_palette,io_spritePen_color}; // @[ColorMixer.scala 100:48]
  wire [10:0] _paletteRamAddr_T_16 = {1'h0,io_spritePen_palette,io_spritePen_color[3:0]}; // @[ColorMixer.scala 101:35]
  wire [12:0] _paletteRamAddr_T_19 = {1'h0,io_spritePen_palette,io_spritePen_color[5:0]}; // @[ColorMixer.scala 102:35]
  wire [14:0] _paletteRamAddr_T_21 = 9'h10 == io_gameConfig_granularity ? {{4'd0}, _paletteRamAddr_T_16} :
    _paletteRamAddr_T_13; // @[Mux.scala 81:58]
  wire [14:0] _paletteRamAddr_T_23 = 9'h40 == io_gameConfig_granularity ? {{2'd0}, _paletteRamAddr_T_19} :
    _paletteRamAddr_T_21; // @[Mux.scala 81:58]
  wire [15:0] _paletteRamAddr_T_25 = {io_gameConfig_layer_0_paletteBank,io_layer0Pen_palette,io_layer0Pen_color}; // @[ColorMixer.scala 100:48]
  wire [11:0] _paletteRamAddr_T_28 = {io_gameConfig_layer_0_paletteBank,io_layer0Pen_palette,io_layer0Pen_color[3:0]}; // @[ColorMixer.scala 101:35]
  wire [13:0] _paletteRamAddr_T_31 = {io_gameConfig_layer_0_paletteBank,io_layer0Pen_palette,io_layer0Pen_color[5:0]}; // @[ColorMixer.scala 102:35]
  wire [15:0] _paletteRamAddr_T_33 = 9'h10 == io_gameConfig_granularity ? {{4'd0}, _paletteRamAddr_T_28} :
    _paletteRamAddr_T_25; // @[Mux.scala 81:58]
  wire [15:0] _paletteRamAddr_T_35 = 9'h40 == io_gameConfig_granularity ? {{2'd0}, _paletteRamAddr_T_31} :
    _paletteRamAddr_T_33; // @[Mux.scala 81:58]
  wire [15:0] _paletteRamAddr_T_37 = {io_gameConfig_layer_1_paletteBank,io_layer1Pen_palette,io_layer1Pen_color}; // @[ColorMixer.scala 100:48]
  wire [11:0] _paletteRamAddr_T_40 = {io_gameConfig_layer_1_paletteBank,io_layer1Pen_palette,io_layer1Pen_color[3:0]}; // @[ColorMixer.scala 101:35]
  wire [13:0] _paletteRamAddr_T_43 = {io_gameConfig_layer_1_paletteBank,io_layer1Pen_palette,io_layer1Pen_color[5:0]}; // @[ColorMixer.scala 102:35]
  wire [15:0] _paletteRamAddr_T_45 = 9'h10 == io_gameConfig_granularity ? {{4'd0}, _paletteRamAddr_T_40} :
    _paletteRamAddr_T_37; // @[Mux.scala 81:58]
  wire [15:0] _paletteRamAddr_T_47 = 9'h40 == io_gameConfig_granularity ? {{2'd0}, _paletteRamAddr_T_43} :
    _paletteRamAddr_T_45; // @[Mux.scala 81:58]
  wire [15:0] _paletteRamAddr_T_49 = {io_gameConfig_layer_2_paletteBank,io_layer2Pen_palette,io_layer2Pen_color}; // @[ColorMixer.scala 100:48]
  wire [11:0] _paletteRamAddr_T_52 = {io_gameConfig_layer_2_paletteBank,io_layer2Pen_palette,io_layer2Pen_color[3:0]}; // @[ColorMixer.scala 101:35]
  wire [13:0] _paletteRamAddr_T_55 = {io_gameConfig_layer_2_paletteBank,io_layer2Pen_palette,io_layer2Pen_color[5:0]}; // @[ColorMixer.scala 102:35]
  wire [15:0] _paletteRamAddr_T_57 = 9'h10 == io_gameConfig_granularity ? {{4'd0}, _paletteRamAddr_T_52} :
    _paletteRamAddr_T_49; // @[Mux.scala 81:58]
  wire [15:0] _paletteRamAddr_T_59 = 9'h40 == io_gameConfig_granularity ? {{2'd0}, _paletteRamAddr_T_55} :
    _paletteRamAddr_T_57; // @[Mux.scala 81:58]
  wire [14:0] _paletteRamAddr_T_61 = 4'h0 == index ? _paletteRamAddr_T_11 : 15'h0; // @[Mux.scala 81:58]
  wire [14:0] _paletteRamAddr_T_63 = 4'h1 == index ? _paletteRamAddr_T_23 : _paletteRamAddr_T_61; // @[Mux.scala 81:58]
  wire [15:0] _paletteRamAddr_T_65 = 4'h2 == index ? _paletteRamAddr_T_35 : {{1'd0}, _paletteRamAddr_T_63}; // @[Mux.scala 81:58]
  wire [15:0] _paletteRamAddr_T_67 = 4'h4 == index ? _paletteRamAddr_T_47 : _paletteRamAddr_T_65; // @[Mux.scala 81:58]
  wire [15:0] paletteRamAddr = 4'h8 == index ? _paletteRamAddr_T_59 : _paletteRamAddr_T_67; // @[Mux.scala 81:58]
  reg [15:0] io_dout_REG; // @[ColorMixer.scala 76:21]
  assign io_paletteRam_addr = paletteRamAddr[14:0]; // @[ColorMixer.scala 75:22]
  assign io_dout = io_dout_REG; // @[ColorMixer.scala 76:11]
  always @(posedge clock) begin
    io_dout_REG <= io_paletteRam_dout; // @[ColorMixer.scala 76:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_dout_REG = _RAND_0[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GPU(
  input          clock,
  input          reset,
  input          io_videoClock,
  input          io_layerCtrl_0_enable,
  input  [1:0]   io_layerCtrl_0_format,
  input          io_layerCtrl_0_regs_tileSize,
  input          io_layerCtrl_0_regs_enable,
  input          io_layerCtrl_0_regs_flipX,
  input          io_layerCtrl_0_regs_flipY,
  input          io_layerCtrl_0_regs_rowScrollEnable,
  input          io_layerCtrl_0_regs_rowSelectEnable,
  input  [8:0]   io_layerCtrl_0_regs_scroll_x,
  input  [8:0]   io_layerCtrl_0_regs_scroll_y,
  output [11:0]  io_layerCtrl_0_vram8x8_addr,
  input  [31:0]  io_layerCtrl_0_vram8x8_dout,
  output [9:0]   io_layerCtrl_0_vram16x16_addr,
  input  [31:0]  io_layerCtrl_0_vram16x16_dout,
  output [8:0]   io_layerCtrl_0_lineRam_addr,
  input  [31:0]  io_layerCtrl_0_lineRam_dout,
  output         io_layerCtrl_0_tileRom_rd,
  output [31:0]  io_layerCtrl_0_tileRom_addr,
  input  [63:0]  io_layerCtrl_0_tileRom_dout,
  input          io_layerCtrl_1_enable,
  input  [1:0]   io_layerCtrl_1_format,
  input          io_layerCtrl_1_regs_tileSize,
  input          io_layerCtrl_1_regs_enable,
  input          io_layerCtrl_1_regs_flipX,
  input          io_layerCtrl_1_regs_flipY,
  input          io_layerCtrl_1_regs_rowScrollEnable,
  input          io_layerCtrl_1_regs_rowSelectEnable,
  input  [8:0]   io_layerCtrl_1_regs_scroll_x,
  input  [8:0]   io_layerCtrl_1_regs_scroll_y,
  output [11:0]  io_layerCtrl_1_vram8x8_addr,
  input  [31:0]  io_layerCtrl_1_vram8x8_dout,
  output [9:0]   io_layerCtrl_1_vram16x16_addr,
  input  [31:0]  io_layerCtrl_1_vram16x16_dout,
  output [8:0]   io_layerCtrl_1_lineRam_addr,
  input  [31:0]  io_layerCtrl_1_lineRam_dout,
  output         io_layerCtrl_1_tileRom_rd,
  output [31:0]  io_layerCtrl_1_tileRom_addr,
  input  [63:0]  io_layerCtrl_1_tileRom_dout,
  input          io_layerCtrl_2_enable,
  input  [1:0]   io_layerCtrl_2_format,
  input          io_layerCtrl_2_regs_tileSize,
  input          io_layerCtrl_2_regs_enable,
  input          io_layerCtrl_2_regs_flipX,
  input          io_layerCtrl_2_regs_flipY,
  input          io_layerCtrl_2_regs_rowScrollEnable,
  input          io_layerCtrl_2_regs_rowSelectEnable,
  input  [8:0]   io_layerCtrl_2_regs_scroll_x,
  input  [8:0]   io_layerCtrl_2_regs_scroll_y,
  output [11:0]  io_layerCtrl_2_vram8x8_addr,
  input  [31:0]  io_layerCtrl_2_vram8x8_dout,
  output [9:0]   io_layerCtrl_2_vram16x16_addr,
  input  [31:0]  io_layerCtrl_2_vram16x16_dout,
  output [8:0]   io_layerCtrl_2_lineRam_addr,
  input  [31:0]  io_layerCtrl_2_lineRam_dout,
  output         io_layerCtrl_2_tileRom_rd,
  output [31:0]  io_layerCtrl_2_tileRom_addr,
  input  [63:0]  io_layerCtrl_2_tileRom_dout,
  input          io_spriteCtrl_enable,
  input  [1:0]   io_spriteCtrl_format,
  input          io_spriteCtrl_start,
  input          io_spriteCtrl_zoom,
  input  [8:0]   io_spriteCtrl_regs_offset_x,
  input  [8:0]   io_spriteCtrl_regs_offset_y,
  input  [1:0]   io_spriteCtrl_regs_bank,
  input          io_spriteCtrl_regs_fixed,
  input          io_spriteCtrl_regs_hFlip,
  output         io_spriteCtrl_vram_rd,
  output [11:0]  io_spriteCtrl_vram_addr,
  input  [127:0] io_spriteCtrl_vram_dout,
  output         io_spriteCtrl_tileRom_rd,
  output [31:0]  io_spriteCtrl_tileRom_addr,
  input  [63:0]  io_spriteCtrl_tileRom_dout,
  input          io_spriteCtrl_tileRom_wait_n,
  input          io_spriteCtrl_tileRom_valid,
  output [7:0]   io_spriteCtrl_tileRom_burstLength,
  input          io_spriteCtrl_tileRom_burstDone,
  input  [8:0]   io_gameConfig_granularity,
  input  [1:0]   io_gameConfig_layer_0_paletteBank,
  input  [1:0]   io_gameConfig_layer_1_paletteBank,
  input  [1:0]   io_gameConfig_layer_2_paletteBank,
  input          io_options_rotate,
  input          io_options_flip,
  input          io_video_clockEnable,
  input          io_video_displayEnable,
  input  [8:0]   io_video_pos_x,
  input  [8:0]   io_video_pos_y,
  input          io_video_vBlank,
  input  [8:0]   io_video_regs_size_x,
  input  [8:0]   io_video_regs_size_y,
  output [8:0]   io_spriteLineBuffer_addr,
  input  [15:0]  io_spriteLineBuffer_dout,
  output         io_spriteFrameBuffer_wr,
  output [16:0]  io_spriteFrameBuffer_addr,
  output [15:0]  io_spriteFrameBuffer_din,
  input          io_spriteFrameBuffer_wait_n,
  output         io_systemFrameBuffer_wr,
  output [16:0]  io_systemFrameBuffer_addr,
  output [31:0]  io_systemFrameBuffer_din,
  output [14:0]  io_paletteRam_addr,
  input  [15:0]  io_paletteRam_dout,
  output [23:0]  io_rgb
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  spriteProcessor_clock; // @[GPU.scala 76:31]
  wire  spriteProcessor_reset; // @[GPU.scala 76:31]
  wire  spriteProcessor_io_ctrl_enable; // @[GPU.scala 76:31]
  wire [1:0] spriteProcessor_io_ctrl_format; // @[GPU.scala 76:31]
  wire  spriteProcessor_io_ctrl_start; // @[GPU.scala 76:31]
  wire  spriteProcessor_io_ctrl_zoom; // @[GPU.scala 76:31]
  wire [1:0] spriteProcessor_io_ctrl_regs_bank; // @[GPU.scala 76:31]
  wire  spriteProcessor_io_ctrl_regs_fixed; // @[GPU.scala 76:31]
  wire  spriteProcessor_io_ctrl_regs_hFlip; // @[GPU.scala 76:31]
  wire  spriteProcessor_io_ctrl_vram_rd; // @[GPU.scala 76:31]
  wire [11:0] spriteProcessor_io_ctrl_vram_addr; // @[GPU.scala 76:31]
  wire [127:0] spriteProcessor_io_ctrl_vram_dout; // @[GPU.scala 76:31]
  wire  spriteProcessor_io_ctrl_tileRom_rd; // @[GPU.scala 76:31]
  wire [31:0] spriteProcessor_io_ctrl_tileRom_addr; // @[GPU.scala 76:31]
  wire [63:0] spriteProcessor_io_ctrl_tileRom_dout; // @[GPU.scala 76:31]
  wire  spriteProcessor_io_ctrl_tileRom_wait_n; // @[GPU.scala 76:31]
  wire  spriteProcessor_io_ctrl_tileRom_valid; // @[GPU.scala 76:31]
  wire [7:0] spriteProcessor_io_ctrl_tileRom_burstLength; // @[GPU.scala 76:31]
  wire  spriteProcessor_io_ctrl_tileRom_burstDone; // @[GPU.scala 76:31]
  wire [8:0] spriteProcessor_io_video_regs_size_x; // @[GPU.scala 76:31]
  wire [8:0] spriteProcessor_io_video_regs_size_y; // @[GPU.scala 76:31]
  wire  spriteProcessor_io_frameBuffer_wr; // @[GPU.scala 76:31]
  wire [16:0] spriteProcessor_io_frameBuffer_addr; // @[GPU.scala 76:31]
  wire [15:0] spriteProcessor_io_frameBuffer_din; // @[GPU.scala 76:31]
  wire  spriteProcessor_io_frameBuffer_wait_n; // @[GPU.scala 76:31]
  wire  layerProcessor_0_clock; // @[GPU.scala 84:21]
  wire  layerProcessor_0_io_ctrl_enable; // @[GPU.scala 84:21]
  wire [1:0] layerProcessor_0_io_ctrl_format; // @[GPU.scala 84:21]
  wire  layerProcessor_0_io_ctrl_regs_tileSize; // @[GPU.scala 84:21]
  wire  layerProcessor_0_io_ctrl_regs_enable; // @[GPU.scala 84:21]
  wire  layerProcessor_0_io_ctrl_regs_flipX; // @[GPU.scala 84:21]
  wire  layerProcessor_0_io_ctrl_regs_flipY; // @[GPU.scala 84:21]
  wire  layerProcessor_0_io_ctrl_regs_rowScrollEnable; // @[GPU.scala 84:21]
  wire  layerProcessor_0_io_ctrl_regs_rowSelectEnable; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_0_io_ctrl_regs_scroll_x; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_0_io_ctrl_regs_scroll_y; // @[GPU.scala 84:21]
  wire [11:0] layerProcessor_0_io_ctrl_vram8x8_addr; // @[GPU.scala 84:21]
  wire [31:0] layerProcessor_0_io_ctrl_vram8x8_dout; // @[GPU.scala 84:21]
  wire [9:0] layerProcessor_0_io_ctrl_vram16x16_addr; // @[GPU.scala 84:21]
  wire [31:0] layerProcessor_0_io_ctrl_vram16x16_dout; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_0_io_ctrl_lineRam_addr; // @[GPU.scala 84:21]
  wire [31:0] layerProcessor_0_io_ctrl_lineRam_dout; // @[GPU.scala 84:21]
  wire  layerProcessor_0_io_ctrl_tileRom_rd; // @[GPU.scala 84:21]
  wire [31:0] layerProcessor_0_io_ctrl_tileRom_addr; // @[GPU.scala 84:21]
  wire [63:0] layerProcessor_0_io_ctrl_tileRom_dout; // @[GPU.scala 84:21]
  wire  layerProcessor_0_io_video_clockEnable; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_0_io_video_pos_x; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_0_io_video_pos_y; // @[GPU.scala 84:21]
  wire  layerProcessor_0_io_video_vBlank; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_0_io_video_regs_size_x; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_0_io_video_regs_size_y; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_0_io_spriteOffset_x; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_0_io_spriteOffset_y; // @[GPU.scala 84:21]
  wire [1:0] layerProcessor_0_io_pen_priority; // @[GPU.scala 84:21]
  wire [5:0] layerProcessor_0_io_pen_palette; // @[GPU.scala 84:21]
  wire [7:0] layerProcessor_0_io_pen_color; // @[GPU.scala 84:21]
  wire  layerProcessor_1_clock; // @[GPU.scala 84:21]
  wire  layerProcessor_1_io_ctrl_enable; // @[GPU.scala 84:21]
  wire [1:0] layerProcessor_1_io_ctrl_format; // @[GPU.scala 84:21]
  wire  layerProcessor_1_io_ctrl_regs_tileSize; // @[GPU.scala 84:21]
  wire  layerProcessor_1_io_ctrl_regs_enable; // @[GPU.scala 84:21]
  wire  layerProcessor_1_io_ctrl_regs_flipX; // @[GPU.scala 84:21]
  wire  layerProcessor_1_io_ctrl_regs_flipY; // @[GPU.scala 84:21]
  wire  layerProcessor_1_io_ctrl_regs_rowScrollEnable; // @[GPU.scala 84:21]
  wire  layerProcessor_1_io_ctrl_regs_rowSelectEnable; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_1_io_ctrl_regs_scroll_x; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_1_io_ctrl_regs_scroll_y; // @[GPU.scala 84:21]
  wire [11:0] layerProcessor_1_io_ctrl_vram8x8_addr; // @[GPU.scala 84:21]
  wire [31:0] layerProcessor_1_io_ctrl_vram8x8_dout; // @[GPU.scala 84:21]
  wire [9:0] layerProcessor_1_io_ctrl_vram16x16_addr; // @[GPU.scala 84:21]
  wire [31:0] layerProcessor_1_io_ctrl_vram16x16_dout; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_1_io_ctrl_lineRam_addr; // @[GPU.scala 84:21]
  wire [31:0] layerProcessor_1_io_ctrl_lineRam_dout; // @[GPU.scala 84:21]
  wire  layerProcessor_1_io_ctrl_tileRom_rd; // @[GPU.scala 84:21]
  wire [31:0] layerProcessor_1_io_ctrl_tileRom_addr; // @[GPU.scala 84:21]
  wire [63:0] layerProcessor_1_io_ctrl_tileRom_dout; // @[GPU.scala 84:21]
  wire  layerProcessor_1_io_video_clockEnable; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_1_io_video_pos_x; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_1_io_video_pos_y; // @[GPU.scala 84:21]
  wire  layerProcessor_1_io_video_vBlank; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_1_io_video_regs_size_x; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_1_io_video_regs_size_y; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_1_io_spriteOffset_x; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_1_io_spriteOffset_y; // @[GPU.scala 84:21]
  wire [1:0] layerProcessor_1_io_pen_priority; // @[GPU.scala 84:21]
  wire [5:0] layerProcessor_1_io_pen_palette; // @[GPU.scala 84:21]
  wire [7:0] layerProcessor_1_io_pen_color; // @[GPU.scala 84:21]
  wire  layerProcessor_2_clock; // @[GPU.scala 84:21]
  wire  layerProcessor_2_io_ctrl_enable; // @[GPU.scala 84:21]
  wire [1:0] layerProcessor_2_io_ctrl_format; // @[GPU.scala 84:21]
  wire  layerProcessor_2_io_ctrl_regs_tileSize; // @[GPU.scala 84:21]
  wire  layerProcessor_2_io_ctrl_regs_enable; // @[GPU.scala 84:21]
  wire  layerProcessor_2_io_ctrl_regs_flipX; // @[GPU.scala 84:21]
  wire  layerProcessor_2_io_ctrl_regs_flipY; // @[GPU.scala 84:21]
  wire  layerProcessor_2_io_ctrl_regs_rowScrollEnable; // @[GPU.scala 84:21]
  wire  layerProcessor_2_io_ctrl_regs_rowSelectEnable; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_2_io_ctrl_regs_scroll_x; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_2_io_ctrl_regs_scroll_y; // @[GPU.scala 84:21]
  wire [11:0] layerProcessor_2_io_ctrl_vram8x8_addr; // @[GPU.scala 84:21]
  wire [31:0] layerProcessor_2_io_ctrl_vram8x8_dout; // @[GPU.scala 84:21]
  wire [9:0] layerProcessor_2_io_ctrl_vram16x16_addr; // @[GPU.scala 84:21]
  wire [31:0] layerProcessor_2_io_ctrl_vram16x16_dout; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_2_io_ctrl_lineRam_addr; // @[GPU.scala 84:21]
  wire [31:0] layerProcessor_2_io_ctrl_lineRam_dout; // @[GPU.scala 84:21]
  wire  layerProcessor_2_io_ctrl_tileRom_rd; // @[GPU.scala 84:21]
  wire [31:0] layerProcessor_2_io_ctrl_tileRom_addr; // @[GPU.scala 84:21]
  wire [63:0] layerProcessor_2_io_ctrl_tileRom_dout; // @[GPU.scala 84:21]
  wire  layerProcessor_2_io_video_clockEnable; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_2_io_video_pos_x; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_2_io_video_pos_y; // @[GPU.scala 84:21]
  wire  layerProcessor_2_io_video_vBlank; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_2_io_video_regs_size_x; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_2_io_video_regs_size_y; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_2_io_spriteOffset_x; // @[GPU.scala 84:21]
  wire [8:0] layerProcessor_2_io_spriteOffset_y; // @[GPU.scala 84:21]
  wire [1:0] layerProcessor_2_io_pen_priority; // @[GPU.scala 84:21]
  wire [5:0] layerProcessor_2_io_pen_palette; // @[GPU.scala 84:21]
  wire [7:0] layerProcessor_2_io_pen_color; // @[GPU.scala 84:21]
  wire  colorMixer_clock; // @[GPU.scala 92:28]
  wire [8:0] colorMixer_io_gameConfig_granularity; // @[GPU.scala 92:28]
  wire [1:0] colorMixer_io_gameConfig_layer_0_paletteBank; // @[GPU.scala 92:28]
  wire [1:0] colorMixer_io_gameConfig_layer_1_paletteBank; // @[GPU.scala 92:28]
  wire [1:0] colorMixer_io_gameConfig_layer_2_paletteBank; // @[GPU.scala 92:28]
  wire [1:0] colorMixer_io_spritePen_priority; // @[GPU.scala 92:28]
  wire [5:0] colorMixer_io_spritePen_palette; // @[GPU.scala 92:28]
  wire [7:0] colorMixer_io_spritePen_color; // @[GPU.scala 92:28]
  wire [1:0] colorMixer_io_layer0Pen_priority; // @[GPU.scala 92:28]
  wire [5:0] colorMixer_io_layer0Pen_palette; // @[GPU.scala 92:28]
  wire [7:0] colorMixer_io_layer0Pen_color; // @[GPU.scala 92:28]
  wire [1:0] colorMixer_io_layer1Pen_priority; // @[GPU.scala 92:28]
  wire [5:0] colorMixer_io_layer1Pen_palette; // @[GPU.scala 92:28]
  wire [7:0] colorMixer_io_layer1Pen_color; // @[GPU.scala 92:28]
  wire [1:0] colorMixer_io_layer2Pen_priority; // @[GPU.scala 92:28]
  wire [5:0] colorMixer_io_layer2Pen_palette; // @[GPU.scala 92:28]
  wire [7:0] colorMixer_io_layer2Pen_color; // @[GPU.scala 92:28]
  wire [14:0] colorMixer_io_paletteRam_addr; // @[GPU.scala 92:28]
  wire [15:0] colorMixer_io_paletteRam_dout; // @[GPU.scala 92:28]
  wire [15:0] colorMixer_io_dout; // @[GPU.scala 92:28]
  reg  io_systemFrameBuffer_wr_REG; // @[GPU.scala 105:39]
  wire [8:0] _io_systemFrameBuffer_addr_x__T_1 = io_video_regs_size_x - io_video_pos_x; // @[GPU.scala 129:21]
  wire [8:0] io_systemFrameBuffer_addr_x_ = _io_systemFrameBuffer_addr_x__T_1 - 9'h1; // @[GPU.scala 129:29]
  wire [8:0] _io_systemFrameBuffer_addr_y__T_1 = io_video_regs_size_y - io_video_pos_y; // @[GPU.scala 130:21]
  wire [8:0] io_systemFrameBuffer_addr_y_ = _io_systemFrameBuffer_addr_y__T_1 - 9'h1; // @[GPU.scala 130:29]
  wire [17:0] _io_systemFrameBuffer_addr_T = io_video_pos_x * io_video_regs_size_y; // @[GPU.scala 132:20]
  wire [17:0] _GEN_0 = {{9'd0}, io_systemFrameBuffer_addr_y_}; // @[GPU.scala 132:30]
  wire [17:0] _io_systemFrameBuffer_addr_T_2 = _io_systemFrameBuffer_addr_T + _GEN_0; // @[GPU.scala 132:30]
  wire [17:0] _io_systemFrameBuffer_addr_T_3 = io_systemFrameBuffer_addr_x_ * io_video_regs_size_y; // @[GPU.scala 132:40]
  wire [17:0] _GEN_1 = {{9'd0}, io_video_pos_y}; // @[GPU.scala 132:50]
  wire [17:0] _io_systemFrameBuffer_addr_T_5 = _io_systemFrameBuffer_addr_T_3 + _GEN_1; // @[GPU.scala 132:50]
  wire [17:0] _io_systemFrameBuffer_addr_T_7 = io_systemFrameBuffer_addr_y_ * io_video_regs_size_x; // @[GPU.scala 133:21]
  wire [17:0] _GEN_2 = {{9'd0}, io_systemFrameBuffer_addr_x_}; // @[GPU.scala 133:31]
  wire [17:0] _io_systemFrameBuffer_addr_T_9 = _io_systemFrameBuffer_addr_T_7 + _GEN_2; // @[GPU.scala 133:31]
  wire [17:0] _io_systemFrameBuffer_addr_T_10 = io_video_pos_y * io_video_regs_size_x; // @[GPU.scala 133:40]
  wire [17:0] _GEN_3 = {{9'd0}, io_video_pos_x}; // @[GPU.scala 133:50]
  wire [17:0] _io_systemFrameBuffer_addr_T_12 = _io_systemFrameBuffer_addr_T_10 + _GEN_3; // @[GPU.scala 133:50]
  reg [17:0] io_systemFrameBuffer_addr_REG; // @[GPU.scala 106:41]
  wire [7:0] io_systemFrameBuffer_din_b = {colorMixer_io_dout[4:0],colorMixer_io_dout[4:2]}; // @[GPU.scala 157:24]
  wire [23:0] _io_systemFrameBuffer_din_T = {colorMixer_io_dout[4:0],colorMixer_io_dout[4:2],colorMixer_io_dout[14:10],
    colorMixer_io_dout[14:12],colorMixer_io_dout[9:5],colorMixer_io_dout[9:7]}; // @[Cat.scala 33:92]
  reg [31:0] io_systemFrameBuffer_din_REG; // @[GPU.scala 108:40]
  wire [15:0] _io_rgb_T = {colorMixer_io_dout[9:5],colorMixer_io_dout[9:7],colorMixer_io_dout[14:10],colorMixer_io_dout[
    14:12]}; // @[GPU.scala 147:7]
  SpriteProcessor spriteProcessor ( // @[GPU.scala 76:31]
    .clock(spriteProcessor_clock),
    .reset(spriteProcessor_reset),
    .io_ctrl_enable(spriteProcessor_io_ctrl_enable),
    .io_ctrl_format(spriteProcessor_io_ctrl_format),
    .io_ctrl_start(spriteProcessor_io_ctrl_start),
    .io_ctrl_zoom(spriteProcessor_io_ctrl_zoom),
    .io_ctrl_regs_bank(spriteProcessor_io_ctrl_regs_bank),
    .io_ctrl_regs_fixed(spriteProcessor_io_ctrl_regs_fixed),
    .io_ctrl_regs_hFlip(spriteProcessor_io_ctrl_regs_hFlip),
    .io_ctrl_vram_rd(spriteProcessor_io_ctrl_vram_rd),
    .io_ctrl_vram_addr(spriteProcessor_io_ctrl_vram_addr),
    .io_ctrl_vram_dout(spriteProcessor_io_ctrl_vram_dout),
    .io_ctrl_tileRom_rd(spriteProcessor_io_ctrl_tileRom_rd),
    .io_ctrl_tileRom_addr(spriteProcessor_io_ctrl_tileRom_addr),
    .io_ctrl_tileRom_dout(spriteProcessor_io_ctrl_tileRom_dout),
    .io_ctrl_tileRom_wait_n(spriteProcessor_io_ctrl_tileRom_wait_n),
    .io_ctrl_tileRom_valid(spriteProcessor_io_ctrl_tileRom_valid),
    .io_ctrl_tileRom_burstLength(spriteProcessor_io_ctrl_tileRom_burstLength),
    .io_ctrl_tileRom_burstDone(spriteProcessor_io_ctrl_tileRom_burstDone),
    .io_video_regs_size_x(spriteProcessor_io_video_regs_size_x),
    .io_video_regs_size_y(spriteProcessor_io_video_regs_size_y),
    .io_frameBuffer_wr(spriteProcessor_io_frameBuffer_wr),
    .io_frameBuffer_addr(spriteProcessor_io_frameBuffer_addr),
    .io_frameBuffer_din(spriteProcessor_io_frameBuffer_din),
    .io_frameBuffer_wait_n(spriteProcessor_io_frameBuffer_wait_n)
  );
  LayerProcessor layerProcessor_0 ( // @[GPU.scala 84:21]
    .clock(layerProcessor_0_clock),
    .io_ctrl_enable(layerProcessor_0_io_ctrl_enable),
    .io_ctrl_format(layerProcessor_0_io_ctrl_format),
    .io_ctrl_regs_tileSize(layerProcessor_0_io_ctrl_regs_tileSize),
    .io_ctrl_regs_enable(layerProcessor_0_io_ctrl_regs_enable),
    .io_ctrl_regs_flipX(layerProcessor_0_io_ctrl_regs_flipX),
    .io_ctrl_regs_flipY(layerProcessor_0_io_ctrl_regs_flipY),
    .io_ctrl_regs_rowScrollEnable(layerProcessor_0_io_ctrl_regs_rowScrollEnable),
    .io_ctrl_regs_rowSelectEnable(layerProcessor_0_io_ctrl_regs_rowSelectEnable),
    .io_ctrl_regs_scroll_x(layerProcessor_0_io_ctrl_regs_scroll_x),
    .io_ctrl_regs_scroll_y(layerProcessor_0_io_ctrl_regs_scroll_y),
    .io_ctrl_vram8x8_addr(layerProcessor_0_io_ctrl_vram8x8_addr),
    .io_ctrl_vram8x8_dout(layerProcessor_0_io_ctrl_vram8x8_dout),
    .io_ctrl_vram16x16_addr(layerProcessor_0_io_ctrl_vram16x16_addr),
    .io_ctrl_vram16x16_dout(layerProcessor_0_io_ctrl_vram16x16_dout),
    .io_ctrl_lineRam_addr(layerProcessor_0_io_ctrl_lineRam_addr),
    .io_ctrl_lineRam_dout(layerProcessor_0_io_ctrl_lineRam_dout),
    .io_ctrl_tileRom_rd(layerProcessor_0_io_ctrl_tileRom_rd),
    .io_ctrl_tileRom_addr(layerProcessor_0_io_ctrl_tileRom_addr),
    .io_ctrl_tileRom_dout(layerProcessor_0_io_ctrl_tileRom_dout),
    .io_video_clockEnable(layerProcessor_0_io_video_clockEnable),
    .io_video_pos_x(layerProcessor_0_io_video_pos_x),
    .io_video_pos_y(layerProcessor_0_io_video_pos_y),
    .io_video_vBlank(layerProcessor_0_io_video_vBlank),
    .io_video_regs_size_x(layerProcessor_0_io_video_regs_size_x),
    .io_video_regs_size_y(layerProcessor_0_io_video_regs_size_y),
    .io_spriteOffset_x(layerProcessor_0_io_spriteOffset_x),
    .io_spriteOffset_y(layerProcessor_0_io_spriteOffset_y),
    .io_pen_priority(layerProcessor_0_io_pen_priority),
    .io_pen_palette(layerProcessor_0_io_pen_palette),
    .io_pen_color(layerProcessor_0_io_pen_color)
  );
  LayerProcessor_1 layerProcessor_1 ( // @[GPU.scala 84:21]
    .clock(layerProcessor_1_clock),
    .io_ctrl_enable(layerProcessor_1_io_ctrl_enable),
    .io_ctrl_format(layerProcessor_1_io_ctrl_format),
    .io_ctrl_regs_tileSize(layerProcessor_1_io_ctrl_regs_tileSize),
    .io_ctrl_regs_enable(layerProcessor_1_io_ctrl_regs_enable),
    .io_ctrl_regs_flipX(layerProcessor_1_io_ctrl_regs_flipX),
    .io_ctrl_regs_flipY(layerProcessor_1_io_ctrl_regs_flipY),
    .io_ctrl_regs_rowScrollEnable(layerProcessor_1_io_ctrl_regs_rowScrollEnable),
    .io_ctrl_regs_rowSelectEnable(layerProcessor_1_io_ctrl_regs_rowSelectEnable),
    .io_ctrl_regs_scroll_x(layerProcessor_1_io_ctrl_regs_scroll_x),
    .io_ctrl_regs_scroll_y(layerProcessor_1_io_ctrl_regs_scroll_y),
    .io_ctrl_vram8x8_addr(layerProcessor_1_io_ctrl_vram8x8_addr),
    .io_ctrl_vram8x8_dout(layerProcessor_1_io_ctrl_vram8x8_dout),
    .io_ctrl_vram16x16_addr(layerProcessor_1_io_ctrl_vram16x16_addr),
    .io_ctrl_vram16x16_dout(layerProcessor_1_io_ctrl_vram16x16_dout),
    .io_ctrl_lineRam_addr(layerProcessor_1_io_ctrl_lineRam_addr),
    .io_ctrl_lineRam_dout(layerProcessor_1_io_ctrl_lineRam_dout),
    .io_ctrl_tileRom_rd(layerProcessor_1_io_ctrl_tileRom_rd),
    .io_ctrl_tileRom_addr(layerProcessor_1_io_ctrl_tileRom_addr),
    .io_ctrl_tileRom_dout(layerProcessor_1_io_ctrl_tileRom_dout),
    .io_video_clockEnable(layerProcessor_1_io_video_clockEnable),
    .io_video_pos_x(layerProcessor_1_io_video_pos_x),
    .io_video_pos_y(layerProcessor_1_io_video_pos_y),
    .io_video_vBlank(layerProcessor_1_io_video_vBlank),
    .io_video_regs_size_x(layerProcessor_1_io_video_regs_size_x),
    .io_video_regs_size_y(layerProcessor_1_io_video_regs_size_y),
    .io_spriteOffset_x(layerProcessor_1_io_spriteOffset_x),
    .io_spriteOffset_y(layerProcessor_1_io_spriteOffset_y),
    .io_pen_priority(layerProcessor_1_io_pen_priority),
    .io_pen_palette(layerProcessor_1_io_pen_palette),
    .io_pen_color(layerProcessor_1_io_pen_color)
  );
  LayerProcessor_2 layerProcessor_2 ( // @[GPU.scala 84:21]
    .clock(layerProcessor_2_clock),
    .io_ctrl_enable(layerProcessor_2_io_ctrl_enable),
    .io_ctrl_format(layerProcessor_2_io_ctrl_format),
    .io_ctrl_regs_tileSize(layerProcessor_2_io_ctrl_regs_tileSize),
    .io_ctrl_regs_enable(layerProcessor_2_io_ctrl_regs_enable),
    .io_ctrl_regs_flipX(layerProcessor_2_io_ctrl_regs_flipX),
    .io_ctrl_regs_flipY(layerProcessor_2_io_ctrl_regs_flipY),
    .io_ctrl_regs_rowScrollEnable(layerProcessor_2_io_ctrl_regs_rowScrollEnable),
    .io_ctrl_regs_rowSelectEnable(layerProcessor_2_io_ctrl_regs_rowSelectEnable),
    .io_ctrl_regs_scroll_x(layerProcessor_2_io_ctrl_regs_scroll_x),
    .io_ctrl_regs_scroll_y(layerProcessor_2_io_ctrl_regs_scroll_y),
    .io_ctrl_vram8x8_addr(layerProcessor_2_io_ctrl_vram8x8_addr),
    .io_ctrl_vram8x8_dout(layerProcessor_2_io_ctrl_vram8x8_dout),
    .io_ctrl_vram16x16_addr(layerProcessor_2_io_ctrl_vram16x16_addr),
    .io_ctrl_vram16x16_dout(layerProcessor_2_io_ctrl_vram16x16_dout),
    .io_ctrl_lineRam_addr(layerProcessor_2_io_ctrl_lineRam_addr),
    .io_ctrl_lineRam_dout(layerProcessor_2_io_ctrl_lineRam_dout),
    .io_ctrl_tileRom_rd(layerProcessor_2_io_ctrl_tileRom_rd),
    .io_ctrl_tileRom_addr(layerProcessor_2_io_ctrl_tileRom_addr),
    .io_ctrl_tileRom_dout(layerProcessor_2_io_ctrl_tileRom_dout),
    .io_video_clockEnable(layerProcessor_2_io_video_clockEnable),
    .io_video_pos_x(layerProcessor_2_io_video_pos_x),
    .io_video_pos_y(layerProcessor_2_io_video_pos_y),
    .io_video_vBlank(layerProcessor_2_io_video_vBlank),
    .io_video_regs_size_x(layerProcessor_2_io_video_regs_size_x),
    .io_video_regs_size_y(layerProcessor_2_io_video_regs_size_y),
    .io_spriteOffset_x(layerProcessor_2_io_spriteOffset_x),
    .io_spriteOffset_y(layerProcessor_2_io_spriteOffset_y),
    .io_pen_priority(layerProcessor_2_io_pen_priority),
    .io_pen_palette(layerProcessor_2_io_pen_palette),
    .io_pen_color(layerProcessor_2_io_pen_color)
  );
  ColorMixer colorMixer ( // @[GPU.scala 92:28]
    .clock(colorMixer_clock),
    .io_gameConfig_granularity(colorMixer_io_gameConfig_granularity),
    .io_gameConfig_layer_0_paletteBank(colorMixer_io_gameConfig_layer_0_paletteBank),
    .io_gameConfig_layer_1_paletteBank(colorMixer_io_gameConfig_layer_1_paletteBank),
    .io_gameConfig_layer_2_paletteBank(colorMixer_io_gameConfig_layer_2_paletteBank),
    .io_spritePen_priority(colorMixer_io_spritePen_priority),
    .io_spritePen_palette(colorMixer_io_spritePen_palette),
    .io_spritePen_color(colorMixer_io_spritePen_color),
    .io_layer0Pen_priority(colorMixer_io_layer0Pen_priority),
    .io_layer0Pen_palette(colorMixer_io_layer0Pen_palette),
    .io_layer0Pen_color(colorMixer_io_layer0Pen_color),
    .io_layer1Pen_priority(colorMixer_io_layer1Pen_priority),
    .io_layer1Pen_palette(colorMixer_io_layer1Pen_palette),
    .io_layer1Pen_color(colorMixer_io_layer1Pen_color),
    .io_layer2Pen_priority(colorMixer_io_layer2Pen_priority),
    .io_layer2Pen_palette(colorMixer_io_layer2Pen_palette),
    .io_layer2Pen_color(colorMixer_io_layer2Pen_color),
    .io_paletteRam_addr(colorMixer_io_paletteRam_addr),
    .io_paletteRam_dout(colorMixer_io_paletteRam_dout),
    .io_dout(colorMixer_io_dout)
  );
  assign io_layerCtrl_0_vram8x8_addr = layerProcessor_0_io_ctrl_vram8x8_addr; // @[GPU.scala 85:17]
  assign io_layerCtrl_0_vram16x16_addr = layerProcessor_0_io_ctrl_vram16x16_addr; // @[GPU.scala 85:17]
  assign io_layerCtrl_0_lineRam_addr = layerProcessor_0_io_ctrl_lineRam_addr; // @[GPU.scala 85:17]
  assign io_layerCtrl_0_tileRom_rd = layerProcessor_0_io_ctrl_tileRom_rd; // @[GPU.scala 85:17]
  assign io_layerCtrl_0_tileRom_addr = layerProcessor_0_io_ctrl_tileRom_addr; // @[GPU.scala 85:17]
  assign io_layerCtrl_1_vram8x8_addr = layerProcessor_1_io_ctrl_vram8x8_addr; // @[GPU.scala 85:17]
  assign io_layerCtrl_1_vram16x16_addr = layerProcessor_1_io_ctrl_vram16x16_addr; // @[GPU.scala 85:17]
  assign io_layerCtrl_1_lineRam_addr = layerProcessor_1_io_ctrl_lineRam_addr; // @[GPU.scala 85:17]
  assign io_layerCtrl_1_tileRom_rd = layerProcessor_1_io_ctrl_tileRom_rd; // @[GPU.scala 85:17]
  assign io_layerCtrl_1_tileRom_addr = layerProcessor_1_io_ctrl_tileRom_addr; // @[GPU.scala 85:17]
  assign io_layerCtrl_2_vram8x8_addr = layerProcessor_2_io_ctrl_vram8x8_addr; // @[GPU.scala 85:17]
  assign io_layerCtrl_2_vram16x16_addr = layerProcessor_2_io_ctrl_vram16x16_addr; // @[GPU.scala 85:17]
  assign io_layerCtrl_2_lineRam_addr = layerProcessor_2_io_ctrl_lineRam_addr; // @[GPU.scala 85:17]
  assign io_layerCtrl_2_tileRom_rd = layerProcessor_2_io_ctrl_tileRom_rd; // @[GPU.scala 85:17]
  assign io_layerCtrl_2_tileRom_addr = layerProcessor_2_io_ctrl_tileRom_addr; // @[GPU.scala 85:17]
  assign io_spriteCtrl_vram_rd = spriteProcessor_io_ctrl_vram_rd; // @[GPU.scala 77:27]
  assign io_spriteCtrl_vram_addr = spriteProcessor_io_ctrl_vram_addr; // @[GPU.scala 77:27]
  assign io_spriteCtrl_tileRom_rd = spriteProcessor_io_ctrl_tileRom_rd; // @[GPU.scala 77:27]
  assign io_spriteCtrl_tileRom_addr = spriteProcessor_io_ctrl_tileRom_addr; // @[GPU.scala 77:27]
  assign io_spriteCtrl_tileRom_burstLength = spriteProcessor_io_ctrl_tileRom_burstLength; // @[GPU.scala 77:27]
  assign io_spriteLineBuffer_addr = io_video_pos_x; // @[GPU.scala 102:30]
  assign io_spriteFrameBuffer_wr = spriteProcessor_io_frameBuffer_wr; // @[GPU.scala 79:34]
  assign io_spriteFrameBuffer_addr = spriteProcessor_io_frameBuffer_addr; // @[GPU.scala 79:34]
  assign io_spriteFrameBuffer_din = spriteProcessor_io_frameBuffer_din; // @[GPU.scala 79:34]
  assign io_systemFrameBuffer_wr = io_systemFrameBuffer_wr_REG; // @[GPU.scala 105:29]
  assign io_systemFrameBuffer_addr = io_systemFrameBuffer_addr_REG[16:0]; // @[GPU.scala 106:31]
  assign io_systemFrameBuffer_din = io_systemFrameBuffer_din_REG; // @[GPU.scala 108:30]
  assign io_paletteRam_addr = colorMixer_io_paletteRam_addr; // @[GPU.scala 98:30]
  assign io_rgb = {_io_rgb_T,io_systemFrameBuffer_din_b}; // @[GPU.scala 147:12]
  assign spriteProcessor_clock = clock;
  assign spriteProcessor_reset = reset;
  assign spriteProcessor_io_ctrl_enable = io_spriteCtrl_enable; // @[GPU.scala 77:27]
  assign spriteProcessor_io_ctrl_format = io_spriteCtrl_format; // @[GPU.scala 77:27]
  assign spriteProcessor_io_ctrl_start = io_spriteCtrl_start; // @[GPU.scala 77:27]
  assign spriteProcessor_io_ctrl_zoom = io_spriteCtrl_zoom; // @[GPU.scala 77:27]
  assign spriteProcessor_io_ctrl_regs_bank = io_spriteCtrl_regs_bank; // @[GPU.scala 77:27]
  assign spriteProcessor_io_ctrl_regs_fixed = io_spriteCtrl_regs_fixed; // @[GPU.scala 77:27]
  assign spriteProcessor_io_ctrl_regs_hFlip = io_spriteCtrl_regs_hFlip; // @[GPU.scala 77:27]
  assign spriteProcessor_io_ctrl_vram_dout = io_spriteCtrl_vram_dout; // @[GPU.scala 77:27]
  assign spriteProcessor_io_ctrl_tileRom_dout = io_spriteCtrl_tileRom_dout; // @[GPU.scala 77:27]
  assign spriteProcessor_io_ctrl_tileRom_wait_n = io_spriteCtrl_tileRom_wait_n; // @[GPU.scala 77:27]
  assign spriteProcessor_io_ctrl_tileRom_valid = io_spriteCtrl_tileRom_valid; // @[GPU.scala 77:27]
  assign spriteProcessor_io_ctrl_tileRom_burstDone = io_spriteCtrl_tileRom_burstDone; // @[GPU.scala 77:27]
  assign spriteProcessor_io_video_regs_size_x = io_video_regs_size_x; // @[GPU.scala 78:28]
  assign spriteProcessor_io_video_regs_size_y = io_video_regs_size_y; // @[GPU.scala 78:28]
  assign spriteProcessor_io_frameBuffer_wait_n = io_spriteFrameBuffer_wait_n; // @[GPU.scala 79:34]
  assign layerProcessor_0_clock = io_videoClock;
  assign layerProcessor_0_io_ctrl_enable = io_layerCtrl_0_enable; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_format = io_layerCtrl_0_format; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_regs_tileSize = io_layerCtrl_0_regs_tileSize; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_regs_enable = io_layerCtrl_0_regs_enable; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_regs_flipX = io_layerCtrl_0_regs_flipX; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_regs_flipY = io_layerCtrl_0_regs_flipY; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_regs_rowScrollEnable = io_layerCtrl_0_regs_rowScrollEnable; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_regs_rowSelectEnable = io_layerCtrl_0_regs_rowSelectEnable; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_regs_scroll_x = io_layerCtrl_0_regs_scroll_x; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_regs_scroll_y = io_layerCtrl_0_regs_scroll_y; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_vram8x8_dout = io_layerCtrl_0_vram8x8_dout; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_vram16x16_dout = io_layerCtrl_0_vram16x16_dout; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_lineRam_dout = io_layerCtrl_0_lineRam_dout; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_ctrl_tileRom_dout = io_layerCtrl_0_tileRom_dout; // @[GPU.scala 85:17]
  assign layerProcessor_0_io_video_clockEnable = io_video_clockEnable; // @[GPU.scala 86:18]
  assign layerProcessor_0_io_video_pos_x = io_video_pos_x; // @[GPU.scala 86:18]
  assign layerProcessor_0_io_video_pos_y = io_video_pos_y; // @[GPU.scala 86:18]
  assign layerProcessor_0_io_video_vBlank = io_video_vBlank; // @[GPU.scala 86:18]
  assign layerProcessor_0_io_video_regs_size_x = io_video_regs_size_x; // @[GPU.scala 86:18]
  assign layerProcessor_0_io_video_regs_size_y = io_video_regs_size_y; // @[GPU.scala 86:18]
  assign layerProcessor_0_io_spriteOffset_x = io_spriteCtrl_regs_offset_x; // @[GPU.scala 87:25]
  assign layerProcessor_0_io_spriteOffset_y = io_spriteCtrl_regs_offset_y; // @[GPU.scala 87:25]
  assign layerProcessor_1_clock = io_videoClock;
  assign layerProcessor_1_io_ctrl_enable = io_layerCtrl_1_enable; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_format = io_layerCtrl_1_format; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_regs_tileSize = io_layerCtrl_1_regs_tileSize; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_regs_enable = io_layerCtrl_1_regs_enable; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_regs_flipX = io_layerCtrl_1_regs_flipX; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_regs_flipY = io_layerCtrl_1_regs_flipY; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_regs_rowScrollEnable = io_layerCtrl_1_regs_rowScrollEnable; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_regs_rowSelectEnable = io_layerCtrl_1_regs_rowSelectEnable; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_regs_scroll_x = io_layerCtrl_1_regs_scroll_x; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_regs_scroll_y = io_layerCtrl_1_regs_scroll_y; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_vram8x8_dout = io_layerCtrl_1_vram8x8_dout; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_vram16x16_dout = io_layerCtrl_1_vram16x16_dout; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_lineRam_dout = io_layerCtrl_1_lineRam_dout; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_ctrl_tileRom_dout = io_layerCtrl_1_tileRom_dout; // @[GPU.scala 85:17]
  assign layerProcessor_1_io_video_clockEnable = io_video_clockEnable; // @[GPU.scala 86:18]
  assign layerProcessor_1_io_video_pos_x = io_video_pos_x; // @[GPU.scala 86:18]
  assign layerProcessor_1_io_video_pos_y = io_video_pos_y; // @[GPU.scala 86:18]
  assign layerProcessor_1_io_video_vBlank = io_video_vBlank; // @[GPU.scala 86:18]
  assign layerProcessor_1_io_video_regs_size_x = io_video_regs_size_x; // @[GPU.scala 86:18]
  assign layerProcessor_1_io_video_regs_size_y = io_video_regs_size_y; // @[GPU.scala 86:18]
  assign layerProcessor_1_io_spriteOffset_x = io_spriteCtrl_regs_offset_x; // @[GPU.scala 87:25]
  assign layerProcessor_1_io_spriteOffset_y = io_spriteCtrl_regs_offset_y; // @[GPU.scala 87:25]
  assign layerProcessor_2_clock = io_videoClock;
  assign layerProcessor_2_io_ctrl_enable = io_layerCtrl_2_enable; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_format = io_layerCtrl_2_format; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_regs_tileSize = io_layerCtrl_2_regs_tileSize; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_regs_enable = io_layerCtrl_2_regs_enable; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_regs_flipX = io_layerCtrl_2_regs_flipX; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_regs_flipY = io_layerCtrl_2_regs_flipY; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_regs_rowScrollEnable = io_layerCtrl_2_regs_rowScrollEnable; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_regs_rowSelectEnable = io_layerCtrl_2_regs_rowSelectEnable; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_regs_scroll_x = io_layerCtrl_2_regs_scroll_x; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_regs_scroll_y = io_layerCtrl_2_regs_scroll_y; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_vram8x8_dout = io_layerCtrl_2_vram8x8_dout; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_vram16x16_dout = io_layerCtrl_2_vram16x16_dout; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_lineRam_dout = io_layerCtrl_2_lineRam_dout; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_ctrl_tileRom_dout = io_layerCtrl_2_tileRom_dout; // @[GPU.scala 85:17]
  assign layerProcessor_2_io_video_clockEnable = io_video_clockEnable; // @[GPU.scala 86:18]
  assign layerProcessor_2_io_video_pos_x = io_video_pos_x; // @[GPU.scala 86:18]
  assign layerProcessor_2_io_video_pos_y = io_video_pos_y; // @[GPU.scala 86:18]
  assign layerProcessor_2_io_video_vBlank = io_video_vBlank; // @[GPU.scala 86:18]
  assign layerProcessor_2_io_video_regs_size_x = io_video_regs_size_x; // @[GPU.scala 86:18]
  assign layerProcessor_2_io_video_regs_size_y = io_video_regs_size_y; // @[GPU.scala 86:18]
  assign layerProcessor_2_io_spriteOffset_x = io_spriteCtrl_regs_offset_x; // @[GPU.scala 87:25]
  assign layerProcessor_2_io_spriteOffset_y = io_spriteCtrl_regs_offset_y; // @[GPU.scala 87:25]
  assign colorMixer_clock = io_videoClock;
  assign colorMixer_io_gameConfig_granularity = io_gameConfig_granularity; // @[GPU.scala 93:30]
  assign colorMixer_io_gameConfig_layer_0_paletteBank = io_gameConfig_layer_0_paletteBank; // @[GPU.scala 93:30]
  assign colorMixer_io_gameConfig_layer_1_paletteBank = io_gameConfig_layer_1_paletteBank; // @[GPU.scala 93:30]
  assign colorMixer_io_gameConfig_layer_2_paletteBank = io_gameConfig_layer_2_paletteBank; // @[GPU.scala 93:30]
  assign colorMixer_io_spritePen_priority = io_spriteLineBuffer_dout[15:14]; // @[GPU.scala 94:65]
  assign colorMixer_io_spritePen_palette = io_spriteLineBuffer_dout[13:8]; // @[GPU.scala 94:65]
  assign colorMixer_io_spritePen_color = io_spriteLineBuffer_dout[7:0]; // @[GPU.scala 94:65]
  assign colorMixer_io_layer0Pen_priority = layerProcessor_0_io_pen_priority; // @[GPU.scala 95:29]
  assign colorMixer_io_layer0Pen_palette = layerProcessor_0_io_pen_palette; // @[GPU.scala 95:29]
  assign colorMixer_io_layer0Pen_color = layerProcessor_0_io_pen_color; // @[GPU.scala 95:29]
  assign colorMixer_io_layer1Pen_priority = layerProcessor_1_io_pen_priority; // @[GPU.scala 96:29]
  assign colorMixer_io_layer1Pen_palette = layerProcessor_1_io_pen_palette; // @[GPU.scala 96:29]
  assign colorMixer_io_layer1Pen_color = layerProcessor_1_io_pen_color; // @[GPU.scala 96:29]
  assign colorMixer_io_layer2Pen_priority = layerProcessor_2_io_pen_priority; // @[GPU.scala 97:29]
  assign colorMixer_io_layer2Pen_palette = layerProcessor_2_io_pen_palette; // @[GPU.scala 97:29]
  assign colorMixer_io_layer2Pen_color = layerProcessor_2_io_pen_color; // @[GPU.scala 97:29]
  assign colorMixer_io_paletteRam_dout = io_paletteRam_dout; // @[GPU.scala 98:30]
  always @(posedge io_videoClock) begin
    io_systemFrameBuffer_wr_REG <= io_video_clockEnable & io_video_displayEnable; // @[GPU.scala 105:61]
    if (io_options_rotate) begin // @[GPU.scala 131:8]
      if (io_options_flip) begin // @[GPU.scala 132:10]
        io_systemFrameBuffer_addr_REG <= _io_systemFrameBuffer_addr_T_2;
      end else begin
        io_systemFrameBuffer_addr_REG <= _io_systemFrameBuffer_addr_T_5;
      end
    end else if (io_options_flip) begin // @[GPU.scala 133:10]
      io_systemFrameBuffer_addr_REG <= _io_systemFrameBuffer_addr_T_9;
    end else begin
      io_systemFrameBuffer_addr_REG <= _io_systemFrameBuffer_addr_T_12;
    end
    io_systemFrameBuffer_din_REG <= {{8'd0}, _io_systemFrameBuffer_din_T}; // @[GPU.scala 160:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_systemFrameBuffer_wr_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_systemFrameBuffer_addr_REG = _RAND_1[17:0];
  _RAND_2 = {1{`RANDOM}};
  io_systemFrameBuffer_din_REG = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DualClockFIFO(
  input         clock,
  input         io_readClock,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits
);
  wire [31:0] fifo_data; // @[DualClockFIFO.scala 74:20]
  wire  fifo_rdclk; // @[DualClockFIFO.scala 74:20]
  wire  fifo_rdreq; // @[DualClockFIFO.scala 74:20]
  wire  fifo_wrclk; // @[DualClockFIFO.scala 74:20]
  wire  fifo_wrreq; // @[DualClockFIFO.scala 74:20]
  wire [31:0] fifo_q; // @[DualClockFIFO.scala 74:20]
  wire  fifo_rdempty; // @[DualClockFIFO.scala 74:20]
  wire  fifo_wrfull; // @[DualClockFIFO.scala 74:20]
  dual_clock_fifo #(.DATA_WIDTH(32), .DEPTH(4)) fifo ( // @[DualClockFIFO.scala 74:20]
    .data(fifo_data),
    .rdclk(fifo_rdclk),
    .rdreq(fifo_rdreq),
    .wrclk(fifo_wrclk),
    .wrreq(fifo_wrreq),
    .q(fifo_q),
    .rdempty(fifo_rdempty),
    .wrfull(fifo_wrfull)
  );
  assign io_deq_valid = ~fifo_rdempty; // @[DualClockFIFO.scala 85:19]
  assign io_deq_bits = fifo_q; // @[DualClockFIFO.scala 86:{36,36}]
  assign io_enq_ready = ~fifo_wrfull; // @[DualClockFIFO.scala 79:19]
  assign fifo_data = io_enq_bits; // @[DualClockFIFO.scala 80:16]
  assign fifo_rdclk = io_readClock; // @[DualClockFIFO.scala 83:17]
  assign fifo_rdreq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  assign fifo_wrclk = clock; // @[DualClockFIFO.scala 77:17]
  assign fifo_wrreq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
endmodule
module DualClockFIFO_1(
  input         clock,
  input         io_readClock,
  output        io_deq_valid,
  output [63:0] io_deq_bits,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits
);
  wire [63:0] fifo_data; // @[DualClockFIFO.scala 74:20]
  wire  fifo_rdclk; // @[DualClockFIFO.scala 74:20]
  wire  fifo_rdreq; // @[DualClockFIFO.scala 74:20]
  wire  fifo_wrclk; // @[DualClockFIFO.scala 74:20]
  wire  fifo_wrreq; // @[DualClockFIFO.scala 74:20]
  wire [63:0] fifo_q; // @[DualClockFIFO.scala 74:20]
  wire  fifo_rdempty; // @[DualClockFIFO.scala 74:20]
  wire  fifo_wrfull; // @[DualClockFIFO.scala 74:20]
  dual_clock_fifo #(.DATA_WIDTH(64), .DEPTH(4)) fifo ( // @[DualClockFIFO.scala 74:20]
    .data(fifo_data),
    .rdclk(fifo_rdclk),
    .rdreq(fifo_rdreq),
    .wrclk(fifo_wrclk),
    .wrreq(fifo_wrreq),
    .q(fifo_q),
    .rdempty(fifo_rdempty),
    .wrfull(fifo_wrfull)
  );
  assign io_deq_valid = ~fifo_rdempty; // @[DualClockFIFO.scala 85:19]
  assign io_deq_bits = fifo_q; // @[DualClockFIFO.scala 86:{36,36}]
  assign io_enq_ready = ~fifo_wrfull; // @[DualClockFIFO.scala 79:19]
  assign fifo_data = io_enq_bits; // @[DualClockFIFO.scala 80:16]
  assign fifo_rdclk = io_readClock; // @[DualClockFIFO.scala 83:17]
  assign fifo_rdreq = io_deq_valid; // @[Decoupled.scala 52:35]
  assign fifo_wrclk = clock; // @[DualClockFIFO.scala 77:17]
  assign fifo_wrreq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
endmodule
module Crossing(
  input         clock,
  input         io_targetClock,
  input         io_in_rd,
  input  [31:0] io_in_addr,
  output [63:0] io_in_dout,
  output        io_out_rd,
  output [31:0] io_out_addr,
  input  [63:0] io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid
);
  wire  addrFifo_clock; // @[Crossing.scala 56:52]
  wire  addrFifo_io_readClock; // @[Crossing.scala 56:52]
  wire  addrFifo_io_deq_ready; // @[Crossing.scala 56:52]
  wire  addrFifo_io_deq_valid; // @[Crossing.scala 56:52]
  wire [31:0] addrFifo_io_deq_bits; // @[Crossing.scala 56:52]
  wire  addrFifo_io_enq_ready; // @[Crossing.scala 56:52]
  wire  addrFifo_io_enq_valid; // @[Crossing.scala 56:52]
  wire [31:0] addrFifo_io_enq_bits; // @[Crossing.scala 56:52]
  wire  dataFifo_clock; // @[Crossing.scala 60:43]
  wire  dataFifo_io_readClock; // @[Crossing.scala 60:43]
  wire  dataFifo_io_deq_valid; // @[Crossing.scala 60:43]
  wire [63:0] dataFifo_io_deq_bits; // @[Crossing.scala 60:43]
  wire  dataFifo_io_enq_ready; // @[Crossing.scala 60:43]
  wire  dataFifo_io_enq_valid; // @[Crossing.scala 60:43]
  wire [63:0] dataFifo_io_enq_bits; // @[Crossing.scala 60:43]
  DualClockFIFO addrFifo ( // @[Crossing.scala 56:52]
    .clock(addrFifo_clock),
    .io_readClock(addrFifo_io_readClock),
    .io_deq_ready(addrFifo_io_deq_ready),
    .io_deq_valid(addrFifo_io_deq_valid),
    .io_deq_bits(addrFifo_io_deq_bits),
    .io_enq_ready(addrFifo_io_enq_ready),
    .io_enq_valid(addrFifo_io_enq_valid),
    .io_enq_bits(addrFifo_io_enq_bits)
  );
  DualClockFIFO_1 dataFifo ( // @[Crossing.scala 60:43]
    .clock(dataFifo_clock),
    .io_readClock(dataFifo_io_readClock),
    .io_deq_valid(dataFifo_io_deq_valid),
    .io_deq_bits(dataFifo_io_deq_bits),
    .io_enq_ready(dataFifo_io_enq_ready),
    .io_enq_valid(dataFifo_io_enq_valid),
    .io_enq_bits(dataFifo_io_enq_bits)
  );
  assign io_in_dout = dataFifo_io_deq_bits; // @[Crossing.scala 79:14]
  assign io_out_rd = addrFifo_io_deq_valid; // @[Crossing.scala 69:13]
  assign io_out_addr = addrFifo_io_deq_bits; // @[Crossing.scala 71:15]
  assign addrFifo_clock = io_targetClock;
  assign addrFifo_io_readClock = clock; // @[Crossing.scala 57:25]
  assign addrFifo_io_deq_ready = io_out_wait_n; // @[Crossing.scala 70:25]
  assign addrFifo_io_enq_valid = io_in_rd; // @[Crossing.scala 64:25]
  assign addrFifo_io_enq_bits = io_in_addr; // @[Crossing.scala 66:24]
  assign dataFifo_clock = clock;
  assign dataFifo_io_readClock = io_targetClock; // @[Crossing.scala 61:25]
  assign dataFifo_io_enq_valid = io_out_valid; // @[Crossing.scala 74:25]
  assign dataFifo_io_enq_bits = io_out_dout; // @[Crossing.scala 75:24]
endmodule
module TrueDualPortRam_11(
  input         clock,
  input         io_clockB,
  input         io_portA_wr,
  input  [6:0]  io_portA_addr,
  input  [63:0] io_portA_din,
  input  [8:0]  io_portB_addr,
  output [15:0] io_portB_dout
);
  wire  ram_clk_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_rd_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_wr_a; // @[TrueDualPortRam.scala 99:19]
  wire [6:0] ram_addr_a; // @[TrueDualPortRam.scala 99:19]
  wire [7:0] ram_mask_a; // @[TrueDualPortRam.scala 99:19]
  wire [63:0] ram_din_a; // @[TrueDualPortRam.scala 99:19]
  wire [63:0] ram_dout_a; // @[TrueDualPortRam.scala 99:19]
  wire  ram_clk_b; // @[TrueDualPortRam.scala 99:19]
  wire  ram_rd_b; // @[TrueDualPortRam.scala 99:19]
  wire [8:0] ram_addr_b; // @[TrueDualPortRam.scala 99:19]
  wire [15:0] ram_dout_b; // @[TrueDualPortRam.scala 99:19]
  true_dual_port_ram
    #(.ADDR_WIDTH_A(7), .DEPTH_B(512), .DEPTH_A(128), .DATA_WIDTH_A(64), .DATA_WIDTH_B(16), .MASK_ENABLE("FALSE"), .ADDR_WIDTH_B(9))
    ram ( // @[TrueDualPortRam.scala 99:19]
    .clk_a(ram_clk_a),
    .rd_a(ram_rd_a),
    .wr_a(ram_wr_a),
    .addr_a(ram_addr_a),
    .mask_a(ram_mask_a),
    .din_a(ram_din_a),
    .dout_a(ram_dout_a),
    .clk_b(ram_clk_b),
    .rd_b(ram_rd_b),
    .addr_b(ram_addr_b),
    .dout_b(ram_dout_b)
  );
  assign io_portB_dout = ram_dout_b; // @[TrueDualPortRam.scala 110:17]
  assign ram_clk_a = clock; // @[TrueDualPortRam.scala 100:16]
  assign ram_rd_a = 1'h0; // @[TrueDualPortRam.scala 101:15]
  assign ram_wr_a = io_portA_wr; // @[TrueDualPortRam.scala 102:15]
  assign ram_addr_a = io_portA_addr; // @[TrueDualPortRam.scala 103:17]
  assign ram_mask_a = 8'hff; // @[TrueDualPortRam.scala 104:17]
  assign ram_din_a = io_portA_din; // @[TrueDualPortRam.scala 105:16]
  assign ram_clk_b = io_clockB; // @[TrueDualPortRam.scala 107:16]
  assign ram_rd_b = 1'h1; // @[TrueDualPortRam.scala 108:15]
  assign ram_addr_b = io_portB_addr; // @[TrueDualPortRam.scala 109:17]
endmodule
module PageFlipper(
  input         clock,
  input         reset,
  input         io_swapWrite,
  output [31:0] io_addrRead,
  output [31:0] io_addrWrite
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] rdIndexReg; // @[PageFlipper.scala 59:27]
  reg [1:0] wrIndexReg; // @[PageFlipper.scala 60:27]
  wire  _wrIndexReg_T_33 = ~wrIndexReg[0]; // @[PageFlipper.scala 75:21]
  wire [12:0] _io_addrRead_T_1 = {11'h121,rdIndexReg}; // @[PageFlipper.scala 80:37]
  wire [12:0] _io_addrWrite_T_1 = {11'h121,wrIndexReg}; // @[PageFlipper.scala 81:38]
  assign io_addrRead = {_io_addrRead_T_1,19'h0}; // @[PageFlipper.scala 80:57]
  assign io_addrWrite = {_io_addrWrite_T_1,19'h0}; // @[PageFlipper.scala 81:58]
  always @(posedge clock) begin
    if (reset) begin // @[PageFlipper.scala 59:27]
      rdIndexReg <= 2'h0; // @[PageFlipper.scala 59:27]
    end else if (io_swapWrite) begin // @[PageFlipper.scala 73:24]
      rdIndexReg <= {{1'd0}, wrIndexReg[0]}; // @[PageFlipper.scala 74:18]
    end
    if (reset) begin // @[PageFlipper.scala 60:27]
      wrIndexReg <= 2'h1; // @[PageFlipper.scala 60:27]
    end else if (io_swapWrite) begin // @[PageFlipper.scala 73:24]
      wrIndexReg <= {{1'd0}, _wrIndexReg_T_33}; // @[PageFlipper.scala 75:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rdIndexReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  wrIndexReg = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BurstReadDMA_1(
  input         clock,
  input         reset,
  input         io_start,
  output        io_in_rd,
  output [31:0] io_in_addr,
  input  [63:0] io_in_dout,
  input         io_in_wait_n,
  input         io_in_valid,
  input         io_in_burstDone,
  output        io_out_wr,
  output [31:0] io_out_addr,
  output [63:0] io_out_din
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  fifo_clock; // @[BurstReadDMA.scala 69:20]
  wire  fifo_reset; // @[BurstReadDMA.scala 69:20]
  wire  fifo_io_enq_ready; // @[BurstReadDMA.scala 69:20]
  wire  fifo_io_enq_valid; // @[BurstReadDMA.scala 69:20]
  wire [63:0] fifo_io_enq_bits; // @[BurstReadDMA.scala 69:20]
  wire  fifo_io_deq_ready; // @[BurstReadDMA.scala 69:20]
  wire  fifo_io_deq_valid; // @[BurstReadDMA.scala 69:20]
  wire [63:0] fifo_io_deq_bits; // @[BurstReadDMA.scala 69:20]
  wire [5:0] fifo_io_count; // @[BurstReadDMA.scala 69:20]
  wire  fifo_io_flush; // @[BurstReadDMA.scala 69:20]
  reg  readEnableReg; // @[BurstReadDMA.scala 62:30]
  reg  writeEnableReg; // @[BurstReadDMA.scala 63:31]
  reg  readPendingReg; // @[BurstReadDMA.scala 64:31]
  wire  fifoAlmostEmpty = fifo_io_count <= 6'h10; // @[BurstReadDMA.scala 70:39]
  wire  busy = readEnableReg | writeEnableReg; // @[BurstReadDMA.scala 73:28]
  wire  start = io_start & ~busy; // @[BurstReadDMA.scala 74:24]
  wire  read = readEnableReg & ~readPendingReg & fifoAlmostEmpty; // @[BurstReadDMA.scala 75:47]
  wire  write = writeEnableReg & fifo_io_deq_valid; // @[BurstReadDMA.scala 76:30]
  wire  effectiveRead = read & io_in_wait_n; // @[BurstReadDMA.scala 77:28]
  reg [6:0] wordCounter; // @[Counter.scala 40:34]
  wire  wrap_wrap = wordCounter == 7'h7f; // @[Counter.scala 45:24]
  wire [6:0] _wrap_value_T_1 = wordCounter + 7'h1; // @[Counter.scala 46:22]
  wire  wordCounterWrap = write & wrap_wrap; // @[Counter.scala 86:{48,55}]
  reg [2:0] burstCounter; // @[Counter.scala 40:34]
  wire  wrap_wrap_1 = burstCounter == 3'h7; // @[Counter.scala 45:24]
  wire [2:0] _wrap_value_T_3 = burstCounter + 3'h1; // @[Counter.scala 46:22]
  wire  burstCounterWrap = io_in_burstDone & wrap_wrap_1; // @[Counter.scala 86:{48,55}]
  wire [9:0] readAddr = {burstCounter, 7'h0}; // @[BurstReadDMA.scala 87:19]
  wire [9:0] writeAddr = {wordCounter, 3'h0}; // @[BurstReadDMA.scala 93:18]
  wire  _GEN_8 = burstCounterWrap ? 1'h0 : readEnableReg; // @[BurstReadDMA.scala 100:{70,86} 62:30]
  wire  _GEN_9 = start | _GEN_8; // @[BurstReadDMA.scala 100:{15,31}]
  wire  _GEN_10 = wordCounterWrap ? 1'h0 : writeEnableReg; // @[BurstReadDMA.scala 101:{70,87} 63:31]
  wire  _GEN_11 = start | _GEN_10; // @[BurstReadDMA.scala 101:{15,32}]
  wire  _GEN_12 = effectiveRead | readPendingReg; // @[BurstReadDMA.scala 106:29 107:20 64:31]
  Queue fifo ( // @[BurstReadDMA.scala 69:20]
    .clock(fifo_clock),
    .reset(fifo_reset),
    .io_enq_ready(fifo_io_enq_ready),
    .io_enq_valid(fifo_io_enq_valid),
    .io_enq_bits(fifo_io_enq_bits),
    .io_deq_ready(fifo_io_deq_ready),
    .io_deq_valid(fifo_io_deq_valid),
    .io_deq_bits(fifo_io_deq_bits),
    .io_count(fifo_io_count),
    .io_flush(fifo_io_flush)
  );
  assign io_in_rd = readEnableReg & ~readPendingReg & fifoAlmostEmpty; // @[BurstReadDMA.scala 75:47]
  assign io_in_addr = {{22'd0}, readAddr}; // @[BurstReadDMA.scala 124:14]
  assign io_out_wr = writeEnableReg & fifo_io_deq_valid; // @[BurstReadDMA.scala 76:30]
  assign io_out_addr = {{22'd0}, writeAddr}; // @[BurstReadDMA.scala 126:15]
  assign io_out_din = fifo_io_deq_bits; // @[BurstReadDMA.scala 127:14]
  assign fifo_clock = clock;
  assign fifo_reset = reset;
  assign fifo_io_enq_valid = io_in_valid & readPendingReg; // @[BurstReadDMA.scala 111:20]
  assign fifo_io_enq_bits = io_in_dout; // @[BurstReadDMA.scala 111:39 Decoupled.scala 66:19]
  assign fifo_io_deq_ready = writeEnableReg & fifo_io_deq_valid; // @[BurstReadDMA.scala 76:30]
  assign fifo_io_flush = io_start & ~busy; // @[BurstReadDMA.scala 74:24]
  always @(posedge clock) begin
    if (reset) begin // @[BurstReadDMA.scala 62:30]
      readEnableReg <= 1'h0; // @[BurstReadDMA.scala 62:30]
    end else begin
      readEnableReg <= _GEN_9;
    end
    if (reset) begin // @[BurstReadDMA.scala 63:31]
      writeEnableReg <= 1'h0; // @[BurstReadDMA.scala 63:31]
    end else begin
      writeEnableReg <= _GEN_11;
    end
    if (reset) begin // @[BurstReadDMA.scala 64:31]
      readPendingReg <= 1'h0; // @[BurstReadDMA.scala 64:31]
    end else if (io_in_burstDone) begin // @[BurstReadDMA.scala 104:25]
      readPendingReg <= 1'h0; // @[BurstReadDMA.scala 105:20]
    end else begin
      readPendingReg <= _GEN_12;
    end
    if (reset) begin // @[Counter.scala 40:34]
      wordCounter <= 7'h0; // @[Counter.scala 40:34]
    end else if (write) begin // @[Counter.scala 86:48]
      wordCounter <= _wrap_value_T_1; // @[Counter.scala 46:13]
    end
    if (reset) begin // @[Counter.scala 40:34]
      burstCounter <= 3'h0; // @[Counter.scala 40:34]
    end else if (io_in_burstDone) begin // @[Counter.scala 86:48]
      burstCounter <= _wrap_value_T_3; // @[Counter.scala 46:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  readEnableReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  writeEnableReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  readPendingReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  wordCounter = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  burstCounter = _RAND_4[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DualClockFIFO_6(
  input         clock,
  input         io_readClock,
  input         io_deq_ready,
  output        io_deq_valid,
  output [16:0] io_deq_bits_addr,
  output [15:0] io_deq_bits_din,
  output [1:0]  io_deq_bits_mask,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_wr,
  input  [16:0] io_enq_bits_addr,
  input  [15:0] io_enq_bits_din
);
  wire [35:0] fifo_data; // @[DualClockFIFO.scala 74:20]
  wire  fifo_rdclk; // @[DualClockFIFO.scala 74:20]
  wire  fifo_rdreq; // @[DualClockFIFO.scala 74:20]
  wire  fifo_wrclk; // @[DualClockFIFO.scala 74:20]
  wire  fifo_wrreq; // @[DualClockFIFO.scala 74:20]
  wire [35:0] fifo_q; // @[DualClockFIFO.scala 74:20]
  wire  fifo_rdempty; // @[DualClockFIFO.scala 74:20]
  wire  fifo_wrfull; // @[DualClockFIFO.scala 74:20]
  wire [17:0] fifo_io_data_lo = {io_enq_bits_din,2'h3}; // @[DualClockFIFO.scala 80:31]
  wire [17:0] fifo_io_data_hi = {io_enq_bits_wr,io_enq_bits_addr}; // @[DualClockFIFO.scala 80:31]
  wire [35:0] _io_deq_bits_WIRE_1 = fifo_q;
  dual_clock_fifo #(.DATA_WIDTH(36), .DEPTH(16)) fifo ( // @[DualClockFIFO.scala 74:20]
    .data(fifo_data),
    .rdclk(fifo_rdclk),
    .rdreq(fifo_rdreq),
    .wrclk(fifo_wrclk),
    .wrreq(fifo_wrreq),
    .q(fifo_q),
    .rdempty(fifo_rdempty),
    .wrfull(fifo_wrfull)
  );
  assign io_deq_valid = ~fifo_rdempty; // @[DualClockFIFO.scala 85:19]
  assign io_deq_bits_addr = _io_deq_bits_WIRE_1[34:18]; // @[DualClockFIFO.scala 86:36]
  assign io_deq_bits_din = _io_deq_bits_WIRE_1[17:2]; // @[DualClockFIFO.scala 86:36]
  assign io_deq_bits_mask = _io_deq_bits_WIRE_1[1:0]; // @[DualClockFIFO.scala 86:36]
  assign io_enq_ready = ~fifo_wrfull; // @[DualClockFIFO.scala 79:19]
  assign fifo_data = {fifo_io_data_hi,fifo_io_data_lo}; // @[DualClockFIFO.scala 80:31]
  assign fifo_rdclk = io_readClock; // @[DualClockFIFO.scala 83:17]
  assign fifo_rdreq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  assign fifo_wrclk = clock; // @[DualClockFIFO.scala 77:17]
  assign fifo_wrreq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
endmodule
module RequestQueue(
  input         clock,
  input         io_enable,
  input         io_readClock,
  input         io_in_wr,
  input  [16:0] io_in_addr,
  input  [15:0] io_in_din,
  output        io_in_wait_n,
  output        io_out_wr,
  output [31:0] io_out_addr,
  output [7:0]  io_out_mask,
  output [63:0] io_out_din,
  input         io_out_wait_n
);
  wire  fifo_clock; // @[RequestQueue.scala 70:20]
  wire  fifo_io_readClock; // @[RequestQueue.scala 70:20]
  wire  fifo_io_deq_ready; // @[RequestQueue.scala 70:20]
  wire  fifo_io_deq_valid; // @[RequestQueue.scala 70:20]
  wire [16:0] fifo_io_deq_bits_addr; // @[RequestQueue.scala 70:20]
  wire [15:0] fifo_io_deq_bits_din; // @[RequestQueue.scala 70:20]
  wire [1:0] fifo_io_deq_bits_mask; // @[RequestQueue.scala 70:20]
  wire  fifo_io_enq_ready; // @[RequestQueue.scala 70:20]
  wire  fifo_io_enq_valid; // @[RequestQueue.scala 70:20]
  wire  fifo_io_enq_bits_wr; // @[RequestQueue.scala 70:20]
  wire [16:0] fifo_io_enq_bits_addr; // @[RequestQueue.scala 70:20]
  wire [15:0] fifo_io_enq_bits_din; // @[RequestQueue.scala 70:20]
  wire [17:0] _io_out_addr_T = {fifo_io_deq_bits_addr, 1'h0}; // @[RequestQueue.scala 83:31]
  wire [31:0] io_out_din_lo = {fifo_io_deq_bits_din,fifo_io_deq_bits_din}; // @[Cat.scala 33:92]
  wire [3:0] _io_out_mask_T_1 = {fifo_io_deq_bits_mask, 2'h0}; // @[RequestQueue.scala 98:28]
  wire [5:0] _io_out_mask_T_2 = {fifo_io_deq_bits_mask, 4'h0}; // @[RequestQueue.scala 99:28]
  wire [7:0] _io_out_mask_T_3 = {fifo_io_deq_bits_mask, 6'h0}; // @[RequestQueue.scala 100:28]
  wire [3:0] _io_out_mask_T_5 = 2'h1 == fifo_io_deq_bits_addr[1:0] ? _io_out_mask_T_1 : {{2'd0}, fifo_io_deq_bits_mask}; // @[Mux.scala 81:58]
  wire [5:0] _io_out_mask_T_7 = 2'h2 == fifo_io_deq_bits_addr[1:0] ? _io_out_mask_T_2 : {{2'd0}, _io_out_mask_T_5}; // @[Mux.scala 81:58]
  DualClockFIFO_6 fifo ( // @[RequestQueue.scala 70:20]
    .clock(fifo_clock),
    .io_readClock(fifo_io_readClock),
    .io_deq_ready(fifo_io_deq_ready),
    .io_deq_valid(fifo_io_deq_valid),
    .io_deq_bits_addr(fifo_io_deq_bits_addr),
    .io_deq_bits_din(fifo_io_deq_bits_din),
    .io_deq_bits_mask(fifo_io_deq_bits_mask),
    .io_enq_ready(fifo_io_enq_ready),
    .io_enq_valid(fifo_io_enq_valid),
    .io_enq_bits_wr(fifo_io_enq_bits_wr),
    .io_enq_bits_addr(fifo_io_enq_bits_addr),
    .io_enq_bits_din(fifo_io_enq_bits_din)
  );
  assign io_in_wait_n = fifo_io_enq_ready; // @[RequestQueue.scala 76:16]
  assign io_out_wr = io_enable & fifo_io_deq_valid; // @[RequestQueue.scala 79:26]
  assign io_out_addr = {{14'd0}, _io_out_addr_T}; // @[RequestQueue.scala 83:15]
  assign io_out_mask = 2'h3 == fifo_io_deq_bits_addr[1:0] ? _io_out_mask_T_3 : {{2'd0}, _io_out_mask_T_7}; // @[Mux.scala 81:58]
  assign io_out_din = {io_out_din_lo,io_out_din_lo}; // @[Cat.scala 33:92]
  assign fifo_clock = clock;
  assign fifo_io_readClock = io_readClock; // @[RequestQueue.scala 71:21]
  assign fifo_io_deq_ready = io_out_wait_n; // @[RequestQueue.scala 80:21]
  assign fifo_io_enq_valid = io_in_wr; // @[RequestQueue.scala 74:21]
  assign fifo_io_enq_bits_wr = io_in_wr; // @[WriteRequest.scala 75:19 76:12]
  assign fifo_io_enq_bits_addr = io_in_addr; // @[WriteRequest.scala 75:19 77:14]
  assign fifo_io_enq_bits_din = io_in_din; // @[WriteRequest.scala 75:19 78:13]
endmodule
module Queue_3(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits,
  output [6:0]  io_count,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:63]; // @[Decoupled.scala 275:44]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:44]
  wire [5:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:44]
  wire [63:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:44]
  wire [63:0] ram_MPORT_data; // @[Decoupled.scala 275:44]
  wire [5:0] ram_MPORT_addr; // @[Decoupled.scala 275:44]
  wire  ram_MPORT_mask; // @[Decoupled.scala 275:44]
  wire  ram_MPORT_en; // @[Decoupled.scala 275:44]
  reg  ram_io_deq_bits_MPORT_en_pipe_0;
  reg [5:0] ram_io_deq_bits_MPORT_addr_pipe_0;
  reg [5:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [5:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 278:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 279:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 280:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 281:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  wire [5:0] _value_T_1 = enq_ptr_value + 6'h1; // @[Counter.scala 77:24]
  wire [5:0] _value_T_3 = deq_ptr_value + 6'h1; // @[Counter.scala 77:24]
  wire [6:0] _deq_ptr_next_T_1 = 7'h40 - 7'h1; // @[Decoupled.scala 308:57]
  wire [6:0] _GEN_15 = {{1'd0}, deq_ptr_value}; // @[Decoupled.scala 308:42]
  wire [5:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 328:32]
  wire [6:0] _io_count_T_1 = maybe_full & ptr_match ? 7'h40 : 7'h0; // @[Decoupled.scala 331:20]
  wire [6:0] _GEN_16 = {{1'd0}, ptr_diff}; // @[Decoupled.scala 331:62]
  assign ram_io_deq_bits_MPORT_en = ram_io_deq_bits_MPORT_en_pipe_0;
  assign ram_io_deq_bits_MPORT_addr = ram_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:44]
  assign ram_MPORT_data = 64'h0;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 305:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 304:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_count = _io_count_T_1 | _GEN_16; // @[Decoupled.scala 331:62]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 275:44]
    end
    ram_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_15 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 308:27]
          ram_io_deq_bits_MPORT_addr_pipe_0 <= 6'h0;
        end else begin
          ram_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_io_deq_bits_MPORT_addr_pipe_0 <= deq_ptr_value;
      end
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 6'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 298:15]
      enq_ptr_value <= 6'h0; // @[Counter.scala 98:11]
    end else if (do_enq) begin // @[Decoupled.scala 288:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 6'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 298:15]
      deq_ptr_value <= 6'h0; // @[Counter.scala 98:11]
    end else if (do_deq) begin // @[Decoupled.scala 292:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 278:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 278:27]
    end else if (io_flush) begin // @[Decoupled.scala 298:15]
      maybe_full <= 1'h0; // @[Decoupled.scala 301:16]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 295:27]
      maybe_full <= do_enq; // @[Decoupled.scala 296:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_io_deq_bits_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_io_deq_bits_MPORT_addr_pipe_0 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BurstWriteDMA(
  input         clock,
  input         reset,
  input         io_start,
  output        io_out_wr,
  output [31:0] io_out_addr,
  output [63:0] io_out_din,
  input         io_out_wait_n,
  input         io_out_burstDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  fifo_clock; // @[BurstWriteDMA.scala 70:20]
  wire  fifo_reset; // @[BurstWriteDMA.scala 70:20]
  wire  fifo_io_enq_ready; // @[BurstWriteDMA.scala 70:20]
  wire  fifo_io_enq_valid; // @[BurstWriteDMA.scala 70:20]
  wire  fifo_io_deq_ready; // @[BurstWriteDMA.scala 70:20]
  wire  fifo_io_deq_valid; // @[BurstWriteDMA.scala 70:20]
  wire [63:0] fifo_io_deq_bits; // @[BurstWriteDMA.scala 70:20]
  wire [6:0] fifo_io_count; // @[BurstWriteDMA.scala 70:20]
  wire  fifo_io_flush; // @[BurstWriteDMA.scala 70:20]
  reg  readEnableReg; // @[BurstWriteDMA.scala 62:30]
  reg  writeEnableReg; // @[BurstWriteDMA.scala 63:31]
  reg  readPendingReg; // @[BurstWriteDMA.scala 64:31]
  reg  writePendingReg; // @[BurstWriteDMA.scala 65:32]
  wire  fifoAlmostFull = fifo_io_count >= 7'h3f; // @[BurstWriteDMA.scala 71:38]
  wire  fifoBurstReady = fifo_io_count == 7'h40; // @[BurstWriteDMA.scala 72:38]
  wire  busy = readEnableReg | writeEnableReg; // @[BurstWriteDMA.scala 75:28]
  wire  start = io_start & ~busy; // @[BurstWriteDMA.scala 76:24]
  wire  read = readEnableReg & (~readPendingReg & fifo_io_enq_ready | ~fifoAlmostFull); // @[BurstWriteDMA.scala 77:28]
  wire  write = writeEnableReg & (writePendingReg | fifoBurstReady); // @[BurstWriteDMA.scala 78:30]
  wire  effectiveWrite = write & io_out_wait_n; // @[BurstWriteDMA.scala 80:30]
  reg [14:0] wordCounter; // @[Counter.scala 40:34]
  wire  wrap_wrap = wordCounter == 15'h7fff; // @[Counter.scala 45:24]
  wire [14:0] _wrap_value_T_1 = wordCounter + 15'h1; // @[Counter.scala 46:22]
  wire  wordCounterWrap = read & wrap_wrap; // @[Counter.scala 86:{48,55}]
  reg [8:0] burstCounter; // @[Counter.scala 40:34]
  wire  wrap_wrap_1 = burstCounter == 9'h1ff; // @[Counter.scala 45:24]
  wire [8:0] _wrap_value_T_3 = burstCounter + 9'h1; // @[Counter.scala 46:22]
  wire  burstCounterWrap = io_out_burstDone & wrap_wrap_1; // @[Counter.scala 86:{48,55}]
  wire [17:0] writeAddr = {burstCounter, 9'h0}; // @[BurstWriteDMA.scala 95:19]
  wire  _GEN_8 = wordCounterWrap ? 1'h0 : readEnableReg; // @[BurstWriteDMA.scala 102:{69,85} 62:30]
  wire  _GEN_9 = start | _GEN_8; // @[BurstWriteDMA.scala 102:{15,31}]
  wire  _GEN_10 = burstCounterWrap ? 1'h0 : writeEnableReg; // @[BurstWriteDMA.scala 103:{71,88} 63:31]
  wire  _GEN_11 = start | _GEN_10; // @[BurstWriteDMA.scala 103:{15,32}]
  wire  _GEN_12 = readPendingReg ? 1'h0 : readPendingReg; // @[BurstWriteDMA.scala 108:45 109:20 64:31]
  wire  _GEN_13 = read | _GEN_12; // @[BurstWriteDMA.scala 106:23 107:20]
  wire  _GEN_14 = effectiveWrite | writePendingReg; // @[BurstWriteDMA.scala 115:30 116:21 65:32]
  Queue_3 fifo ( // @[BurstWriteDMA.scala 70:20]
    .clock(fifo_clock),
    .reset(fifo_reset),
    .io_enq_ready(fifo_io_enq_ready),
    .io_enq_valid(fifo_io_enq_valid),
    .io_deq_ready(fifo_io_deq_ready),
    .io_deq_valid(fifo_io_deq_valid),
    .io_deq_bits(fifo_io_deq_bits),
    .io_count(fifo_io_count),
    .io_flush(fifo_io_flush)
  );
  assign io_out_wr = writeEnableReg & (writePendingReg | fifoBurstReady); // @[BurstWriteDMA.scala 78:30]
  assign io_out_addr = {{14'd0}, writeAddr}; // @[BurstWriteDMA.scala 135:15]
  assign io_out_din = fifo_io_deq_bits; // @[BurstWriteDMA.scala 136:14]
  assign fifo_clock = clock;
  assign fifo_reset = reset;
  assign fifo_io_enq_valid = readPendingReg; // @[BurstWriteDMA.scala 120:20]
  assign fifo_io_deq_ready = write & io_out_wait_n; // @[BurstWriteDMA.scala 80:30]
  assign fifo_io_flush = io_start & ~busy; // @[BurstWriteDMA.scala 76:24]
  always @(posedge clock) begin
    if (reset) begin // @[BurstWriteDMA.scala 62:30]
      readEnableReg <= 1'h0; // @[BurstWriteDMA.scala 62:30]
    end else begin
      readEnableReg <= _GEN_9;
    end
    if (reset) begin // @[BurstWriteDMA.scala 63:31]
      writeEnableReg <= 1'h0; // @[BurstWriteDMA.scala 63:31]
    end else begin
      writeEnableReg <= _GEN_11;
    end
    if (reset) begin // @[BurstWriteDMA.scala 64:31]
      readPendingReg <= 1'h0; // @[BurstWriteDMA.scala 64:31]
    end else begin
      readPendingReg <= _GEN_13;
    end
    if (reset) begin // @[BurstWriteDMA.scala 65:32]
      writePendingReg <= 1'h0; // @[BurstWriteDMA.scala 65:32]
    end else if (io_out_burstDone) begin // @[BurstWriteDMA.scala 113:26]
      writePendingReg <= 1'h0; // @[BurstWriteDMA.scala 114:21]
    end else begin
      writePendingReg <= _GEN_14;
    end
    if (reset) begin // @[Counter.scala 40:34]
      wordCounter <= 15'h0; // @[Counter.scala 40:34]
    end else if (read) begin // @[Counter.scala 86:48]
      wordCounter <= _wrap_value_T_1; // @[Counter.scala 46:13]
    end
    if (reset) begin // @[Counter.scala 40:34]
      burstCounter <= 9'h0; // @[Counter.scala 40:34]
    end else if (io_out_burstDone) begin // @[Counter.scala 86:48]
      burstCounter <= _wrap_value_T_3; // @[Counter.scala 46:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  readEnableReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  writeEnableReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  readPendingReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  writePendingReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wordCounter = _RAND_4[14:0];
  _RAND_5 = {1{`RANDOM}};
  burstCounter = _RAND_5[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BurstMemArbiter_2(
  input         clock,
  input         reset,
  input         io_in_0_rd,
  input  [31:0] io_in_0_addr,
  output [63:0] io_in_0_dout,
  output        io_in_0_wait_n,
  output        io_in_0_valid,
  output        io_in_0_burstDone,
  input         io_in_1_wr,
  input  [31:0] io_in_1_addr,
  input  [63:0] io_in_1_din,
  output        io_in_1_wait_n,
  output        io_in_1_burstDone,
  input         io_in_2_wr,
  input  [31:0] io_in_2_addr,
  input  [7:0]  io_in_2_mask,
  input  [63:0] io_in_2_din,
  output        io_in_2_wait_n,
  output        io_out_rd,
  output        io_out_wr,
  output [31:0] io_out_addr,
  output [7:0]  io_out_mask,
  output [63:0] io_out_din,
  input  [63:0] io_out_dout,
  input         io_out_wait_n,
  input         io_out_valid,
  output [7:0]  io_out_burstLength,
  input         io_out_burstDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  busyReg; // @[BurstMemArbiter.scala 73:24]
  reg [2:0] indexReg; // @[BurstMemArbiter.scala 74:25]
  wire [2:0] _index_enc_T = io_in_2_wr ? 3'h4 : 3'h0; // @[Mux.scala 47:70]
  wire [2:0] _index_enc_T_1 = io_in_1_wr ? 3'h2 : _index_enc_T; // @[Mux.scala 47:70]
  wire [2:0] index_enc = io_in_0_rd ? 3'h1 : _index_enc_T_1; // @[Mux.scala 47:70]
  wire [2:0] index = {index_enc[2],index_enc[1],index_enc[0]}; // @[BurstMemArbiter.scala 77:78]
  wire [2:0] chosen = busyReg ? indexReg : index; // @[BurstMemArbiter.scala 80:19]
  wire  effectiveRequest = ~busyReg & (io_out_rd | io_out_wr) & io_out_wait_n; // @[BurstMemArbiter.scala 83:63]
  wire  _GEN_0 = effectiveRequest | busyReg; // @[BurstMemArbiter.scala 88:32 89:13 73:24]
  wire  io_out_anySelected = chosen[0] | chosen[1] | chosen[2]; // @[BurstMemIO.scala 316:45]
  wire [7:0] _io_out_mem_burstLength_T = chosen[0] ? 8'h10 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_burstLength_T_1 = chosen[1] ? 8'h40 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_burstLength_T_2 = chosen[2] ? 8'h1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_burstLength_T_3 = _io_out_mem_burstLength_T | _io_out_mem_burstLength_T_1; // @[Mux.scala 27:73]
  wire [31:0] _io_out_mem_addr_T = chosen[0] ? io_in_0_addr : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_out_mem_addr_T_1 = chosen[1] ? io_in_1_addr : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_out_mem_addr_T_2 = chosen[2] ? io_in_2_addr : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_out_mem_addr_T_3 = _io_out_mem_addr_T | _io_out_mem_addr_T_1; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_mask_T_1 = chosen[1] ? 8'hff : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _io_out_mem_mask_T_2 = chosen[2] ? io_in_2_mask : 8'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_mem_din_T_1 = chosen[1] ? io_in_1_din : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_out_mem_din_T_2 = chosen[2] ? io_in_2_din : 64'h0; // @[Mux.scala 27:73]
  assign io_in_0_dout = io_out_dout; // @[BurstMemIO.scala 317:19 BurstMemArbiter.scala 96:10]
  assign io_in_0_wait_n = (~io_out_anySelected | chosen[0]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_0_valid = chosen[0] & io_out_valid; // @[BurstMemIO.scala 326:30]
  assign io_in_0_burstDone = chosen[0] & io_out_burstDone; // @[BurstMemIO.scala 327:34]
  assign io_in_1_wait_n = (~io_out_anySelected | chosen[1]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_in_1_burstDone = chosen[1] & io_out_burstDone; // @[BurstMemIO.scala 327:34]
  assign io_in_2_wait_n = (~io_out_anySelected | chosen[2]) & io_out_wait_n; // @[BurstMemIO.scala 325:49]
  assign io_out_rd = chosen[0] & io_in_0_rd; // @[Mux.scala 27:73]
  assign io_out_wr = chosen[1] & io_in_1_wr | chosen[2] & io_in_2_wr; // @[Mux.scala 27:73]
  assign io_out_addr = _io_out_mem_addr_T_3 | _io_out_mem_addr_T_2; // @[Mux.scala 27:73]
  assign io_out_mask = _io_out_mem_mask_T_1 | _io_out_mem_mask_T_2; // @[Mux.scala 27:73]
  assign io_out_din = _io_out_mem_din_T_1 | _io_out_mem_din_T_2; // @[Mux.scala 27:73]
  assign io_out_burstLength = _io_out_mem_burstLength_T_3 | _io_out_mem_burstLength_T_2; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (reset) begin // @[BurstMemArbiter.scala 73:24]
      busyReg <= 1'h0; // @[BurstMemArbiter.scala 73:24]
    end else if (io_out_burstDone) begin // @[BurstMemArbiter.scala 86:26]
      busyReg <= 1'h0; // @[BurstMemArbiter.scala 87:13]
    end else begin
      busyReg <= _GEN_0;
    end
    if (reset) begin // @[BurstMemArbiter.scala 74:25]
      indexReg <= 3'h0; // @[BurstMemArbiter.scala 74:25]
    end else if (!(io_out_burstDone)) begin // @[BurstMemArbiter.scala 86:26]
      if (effectiveRequest) begin // @[BurstMemArbiter.scala 88:32]
        indexReg <= index; // @[BurstMemArbiter.scala 90:14]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busyReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  indexReg = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SpriteFrameBuffer(
  input         clock,
  input         reset,
  input         io_videoClock,
  input         io_enable,
  input         io_swap,
  input  [8:0]  io_video_pos_y,
  input         io_video_hBlank,
  input  [8:0]  io_lineBuffer_addr,
  output [15:0] io_lineBuffer_dout,
  input         io_frameBuffer_wr,
  input  [16:0] io_frameBuffer_addr,
  input  [15:0] io_frameBuffer_din,
  output        io_frameBuffer_wait_n,
  output        io_ddr_rd,
  output        io_ddr_wr,
  output [31:0] io_ddr_addr,
  output [7:0]  io_ddr_mask,
  output [63:0] io_ddr_din,
  input  [63:0] io_ddr_dout,
  input         io_ddr_wait_n,
  input         io_ddr_valid,
  output [7:0]  io_ddr_burstLength,
  input         io_ddr_burstDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  lineBuffer_clock; // @[SpriteFrameBuffer.scala 83:26]
  wire  lineBuffer_io_clockB; // @[SpriteFrameBuffer.scala 83:26]
  wire  lineBuffer_io_portA_wr; // @[SpriteFrameBuffer.scala 83:26]
  wire [6:0] lineBuffer_io_portA_addr; // @[SpriteFrameBuffer.scala 83:26]
  wire [63:0] lineBuffer_io_portA_din; // @[SpriteFrameBuffer.scala 83:26]
  wire [8:0] lineBuffer_io_portB_addr; // @[SpriteFrameBuffer.scala 83:26]
  wire [15:0] lineBuffer_io_portB_dout; // @[SpriteFrameBuffer.scala 83:26]
  wire  pageFlipper_clock; // @[SpriteFrameBuffer.scala 96:27]
  wire  pageFlipper_reset; // @[SpriteFrameBuffer.scala 96:27]
  wire  pageFlipper_io_swapWrite; // @[SpriteFrameBuffer.scala 96:27]
  wire [31:0] pageFlipper_io_addrRead; // @[SpriteFrameBuffer.scala 96:27]
  wire [31:0] pageFlipper_io_addrWrite; // @[SpriteFrameBuffer.scala 96:27]
  wire  lineBufferDma_clock; // @[SpriteFrameBuffer.scala 102:29]
  wire  lineBufferDma_reset; // @[SpriteFrameBuffer.scala 102:29]
  wire  lineBufferDma_io_start; // @[SpriteFrameBuffer.scala 102:29]
  wire  lineBufferDma_io_in_rd; // @[SpriteFrameBuffer.scala 102:29]
  wire [31:0] lineBufferDma_io_in_addr; // @[SpriteFrameBuffer.scala 102:29]
  wire [63:0] lineBufferDma_io_in_dout; // @[SpriteFrameBuffer.scala 102:29]
  wire  lineBufferDma_io_in_wait_n; // @[SpriteFrameBuffer.scala 102:29]
  wire  lineBufferDma_io_in_valid; // @[SpriteFrameBuffer.scala 102:29]
  wire  lineBufferDma_io_in_burstDone; // @[SpriteFrameBuffer.scala 102:29]
  wire  lineBufferDma_io_out_wr; // @[SpriteFrameBuffer.scala 102:29]
  wire [31:0] lineBufferDma_io_out_addr; // @[SpriteFrameBuffer.scala 102:29]
  wire [63:0] lineBufferDma_io_out_din; // @[SpriteFrameBuffer.scala 102:29]
  wire  queue_clock; // @[SpriteFrameBuffer.scala 109:21]
  wire  queue_io_enable; // @[SpriteFrameBuffer.scala 109:21]
  wire  queue_io_readClock; // @[SpriteFrameBuffer.scala 109:21]
  wire  queue_io_in_wr; // @[SpriteFrameBuffer.scala 109:21]
  wire [16:0] queue_io_in_addr; // @[SpriteFrameBuffer.scala 109:21]
  wire [15:0] queue_io_in_din; // @[SpriteFrameBuffer.scala 109:21]
  wire  queue_io_in_wait_n; // @[SpriteFrameBuffer.scala 109:21]
  wire  queue_io_out_wr; // @[SpriteFrameBuffer.scala 109:21]
  wire [31:0] queue_io_out_addr; // @[SpriteFrameBuffer.scala 109:21]
  wire [7:0] queue_io_out_mask; // @[SpriteFrameBuffer.scala 109:21]
  wire [63:0] queue_io_out_din; // @[SpriteFrameBuffer.scala 109:21]
  wire  queue_io_out_wait_n; // @[SpriteFrameBuffer.scala 109:21]
  wire  frameBufferDma_clock; // @[SpriteFrameBuffer.scala 120:30]
  wire  frameBufferDma_reset; // @[SpriteFrameBuffer.scala 120:30]
  wire  frameBufferDma_io_start; // @[SpriteFrameBuffer.scala 120:30]
  wire  frameBufferDma_io_out_wr; // @[SpriteFrameBuffer.scala 120:30]
  wire [31:0] frameBufferDma_io_out_addr; // @[SpriteFrameBuffer.scala 120:30]
  wire [63:0] frameBufferDma_io_out_din; // @[SpriteFrameBuffer.scala 120:30]
  wire  frameBufferDma_io_out_wait_n; // @[SpriteFrameBuffer.scala 120:30]
  wire  frameBufferDma_io_out_burstDone; // @[SpriteFrameBuffer.scala 120:30]
  wire  ddrArbiter_clock; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_reset; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_in_0_rd; // @[SpriteFrameBuffer.scala 130:26]
  wire [31:0] ddrArbiter_io_in_0_addr; // @[SpriteFrameBuffer.scala 130:26]
  wire [63:0] ddrArbiter_io_in_0_dout; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_in_0_wait_n; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_in_0_valid; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_in_0_burstDone; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_in_1_wr; // @[SpriteFrameBuffer.scala 130:26]
  wire [31:0] ddrArbiter_io_in_1_addr; // @[SpriteFrameBuffer.scala 130:26]
  wire [63:0] ddrArbiter_io_in_1_din; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_in_1_wait_n; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_in_1_burstDone; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_in_2_wr; // @[SpriteFrameBuffer.scala 130:26]
  wire [31:0] ddrArbiter_io_in_2_addr; // @[SpriteFrameBuffer.scala 130:26]
  wire [7:0] ddrArbiter_io_in_2_mask; // @[SpriteFrameBuffer.scala 130:26]
  wire [63:0] ddrArbiter_io_in_2_din; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_in_2_wait_n; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_out_rd; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_out_wr; // @[SpriteFrameBuffer.scala 130:26]
  wire [31:0] ddrArbiter_io_out_addr; // @[SpriteFrameBuffer.scala 130:26]
  wire [7:0] ddrArbiter_io_out_mask; // @[SpriteFrameBuffer.scala 130:26]
  wire [63:0] ddrArbiter_io_out_din; // @[SpriteFrameBuffer.scala 130:26]
  wire [63:0] ddrArbiter_io_out_dout; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_out_wait_n; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_out_valid; // @[SpriteFrameBuffer.scala 130:26]
  wire [7:0] ddrArbiter_io_out_burstLength; // @[SpriteFrameBuffer.scala 130:26]
  wire  ddrArbiter_io_out_burstDone; // @[SpriteFrameBuffer.scala 130:26]
  reg  hBlank_r; // @[Reg.scala 19:16]
  reg  hBlank; // @[Reg.scala 19:16]
  reg  hBlankRising_REG; // @[Util.scala 158:44]
  wire  hBlankRising = hBlank & ~hBlankRising_REG; // @[Util.scala 158:33]
  wire [8:0] _lineBufferAddrOffset_T_1 = io_video_pos_y + 9'h1; // @[SpriteFrameBuffer.scala 127:47]
  wire [18:0] lineBufferAddrOffset = {_lineBufferAddrOffset_T_1, 10'h0}; // @[SpriteFrameBuffer.scala 127:54]
  wire [31:0] _mem_T_2 = lineBufferDma_io_in_addr + pageFlipper_io_addrRead; // @[SpriteFrameBuffer.scala 132:35]
  wire [31:0] _GEN_2 = {{13'd0}, lineBufferAddrOffset}; // @[SpriteFrameBuffer.scala 132:61]
  TrueDualPortRam_11 lineBuffer ( // @[SpriteFrameBuffer.scala 83:26]
    .clock(lineBuffer_clock),
    .io_clockB(lineBuffer_io_clockB),
    .io_portA_wr(lineBuffer_io_portA_wr),
    .io_portA_addr(lineBuffer_io_portA_addr),
    .io_portA_din(lineBuffer_io_portA_din),
    .io_portB_addr(lineBuffer_io_portB_addr),
    .io_portB_dout(lineBuffer_io_portB_dout)
  );
  PageFlipper pageFlipper ( // @[SpriteFrameBuffer.scala 96:27]
    .clock(pageFlipper_clock),
    .reset(pageFlipper_reset),
    .io_swapWrite(pageFlipper_io_swapWrite),
    .io_addrRead(pageFlipper_io_addrRead),
    .io_addrWrite(pageFlipper_io_addrWrite)
  );
  BurstReadDMA_1 lineBufferDma ( // @[SpriteFrameBuffer.scala 102:29]
    .clock(lineBufferDma_clock),
    .reset(lineBufferDma_reset),
    .io_start(lineBufferDma_io_start),
    .io_in_rd(lineBufferDma_io_in_rd),
    .io_in_addr(lineBufferDma_io_in_addr),
    .io_in_dout(lineBufferDma_io_in_dout),
    .io_in_wait_n(lineBufferDma_io_in_wait_n),
    .io_in_valid(lineBufferDma_io_in_valid),
    .io_in_burstDone(lineBufferDma_io_in_burstDone),
    .io_out_wr(lineBufferDma_io_out_wr),
    .io_out_addr(lineBufferDma_io_out_addr),
    .io_out_din(lineBufferDma_io_out_din)
  );
  RequestQueue queue ( // @[SpriteFrameBuffer.scala 109:21]
    .clock(queue_clock),
    .io_enable(queue_io_enable),
    .io_readClock(queue_io_readClock),
    .io_in_wr(queue_io_in_wr),
    .io_in_addr(queue_io_in_addr),
    .io_in_din(queue_io_in_din),
    .io_in_wait_n(queue_io_in_wait_n),
    .io_out_wr(queue_io_out_wr),
    .io_out_addr(queue_io_out_addr),
    .io_out_mask(queue_io_out_mask),
    .io_out_din(queue_io_out_din),
    .io_out_wait_n(queue_io_out_wait_n)
  );
  BurstWriteDMA frameBufferDma ( // @[SpriteFrameBuffer.scala 120:30]
    .clock(frameBufferDma_clock),
    .reset(frameBufferDma_reset),
    .io_start(frameBufferDma_io_start),
    .io_out_wr(frameBufferDma_io_out_wr),
    .io_out_addr(frameBufferDma_io_out_addr),
    .io_out_din(frameBufferDma_io_out_din),
    .io_out_wait_n(frameBufferDma_io_out_wait_n),
    .io_out_burstDone(frameBufferDma_io_out_burstDone)
  );
  BurstMemArbiter_2 ddrArbiter ( // @[SpriteFrameBuffer.scala 130:26]
    .clock(ddrArbiter_clock),
    .reset(ddrArbiter_reset),
    .io_in_0_rd(ddrArbiter_io_in_0_rd),
    .io_in_0_addr(ddrArbiter_io_in_0_addr),
    .io_in_0_dout(ddrArbiter_io_in_0_dout),
    .io_in_0_wait_n(ddrArbiter_io_in_0_wait_n),
    .io_in_0_valid(ddrArbiter_io_in_0_valid),
    .io_in_0_burstDone(ddrArbiter_io_in_0_burstDone),
    .io_in_1_wr(ddrArbiter_io_in_1_wr),
    .io_in_1_addr(ddrArbiter_io_in_1_addr),
    .io_in_1_din(ddrArbiter_io_in_1_din),
    .io_in_1_wait_n(ddrArbiter_io_in_1_wait_n),
    .io_in_1_burstDone(ddrArbiter_io_in_1_burstDone),
    .io_in_2_wr(ddrArbiter_io_in_2_wr),
    .io_in_2_addr(ddrArbiter_io_in_2_addr),
    .io_in_2_mask(ddrArbiter_io_in_2_mask),
    .io_in_2_din(ddrArbiter_io_in_2_din),
    .io_in_2_wait_n(ddrArbiter_io_in_2_wait_n),
    .io_out_rd(ddrArbiter_io_out_rd),
    .io_out_wr(ddrArbiter_io_out_wr),
    .io_out_addr(ddrArbiter_io_out_addr),
    .io_out_mask(ddrArbiter_io_out_mask),
    .io_out_din(ddrArbiter_io_out_din),
    .io_out_dout(ddrArbiter_io_out_dout),
    .io_out_wait_n(ddrArbiter_io_out_wait_n),
    .io_out_valid(ddrArbiter_io_out_valid),
    .io_out_burstLength(ddrArbiter_io_out_burstLength),
    .io_out_burstDone(ddrArbiter_io_out_burstDone)
  );
  assign io_lineBuffer_dout = lineBuffer_io_portB_dout; // @[SpriteFrameBuffer.scala 92:23]
  assign io_frameBuffer_wait_n = queue_io_in_wait_n; // @[SpriteFrameBuffer.scala 138:18]
  assign io_ddr_rd = ddrArbiter_io_out_rd; // @[SpriteFrameBuffer.scala 135:5]
  assign io_ddr_wr = ddrArbiter_io_out_wr; // @[SpriteFrameBuffer.scala 135:5]
  assign io_ddr_addr = ddrArbiter_io_out_addr; // @[SpriteFrameBuffer.scala 135:5]
  assign io_ddr_mask = ddrArbiter_io_out_mask; // @[SpriteFrameBuffer.scala 135:5]
  assign io_ddr_din = ddrArbiter_io_out_din; // @[SpriteFrameBuffer.scala 135:5]
  assign io_ddr_burstLength = ddrArbiter_io_out_burstLength; // @[SpriteFrameBuffer.scala 135:5]
  assign lineBuffer_clock = clock;
  assign lineBuffer_io_clockB = io_videoClock; // @[SpriteFrameBuffer.scala 91:24]
  assign lineBuffer_io_portA_wr = lineBufferDma_io_out_wr; // @[AsyncMemIO.scala 236:19 237:12]
  assign lineBuffer_io_portA_addr = lineBufferDma_io_out_addr[9:3]; // @[SpriteFrameBuffer.scala 106:14]
  assign lineBuffer_io_portA_din = lineBufferDma_io_out_din; // @[AsyncMemIO.scala 236:19 241:13]
  assign lineBuffer_io_portB_addr = io_lineBuffer_addr; // @[SpriteFrameBuffer.scala 92:23]
  assign pageFlipper_clock = clock;
  assign pageFlipper_reset = reset;
  assign pageFlipper_io_swapWrite = io_enable & io_swap; // @[SpriteFrameBuffer.scala 99:41]
  assign lineBufferDma_clock = clock;
  assign lineBufferDma_reset = reset;
  assign lineBufferDma_io_start = io_enable & hBlankRising; // @[SpriteFrameBuffer.scala 103:39]
  assign lineBufferDma_io_in_dout = ddrArbiter_io_in_0_dout; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign lineBufferDma_io_in_wait_n = ddrArbiter_io_in_0_wait_n; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign lineBufferDma_io_in_valid = ddrArbiter_io_in_0_valid; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign lineBufferDma_io_in_burstDone = ddrArbiter_io_in_0_burstDone; // @[BurstMemIO.scala 63:19 BurstMemArbiter.scala 68:67]
  assign queue_clock = clock;
  assign queue_io_enable = io_enable; // @[SpriteFrameBuffer.scala 116:19]
  assign queue_io_readClock = clock; // @[SpriteFrameBuffer.scala 117:22]
  assign queue_io_in_wr = io_frameBuffer_wr; // @[SpriteFrameBuffer.scala 138:18]
  assign queue_io_in_addr = io_frameBuffer_addr; // @[SpriteFrameBuffer.scala 138:18]
  assign queue_io_in_din = io_frameBuffer_din; // @[SpriteFrameBuffer.scala 138:18]
  assign queue_io_out_wait_n = ddrArbiter_io_in_2_wait_n; // @[BurstMemIO.scala 156:19 BurstMemArbiter.scala 68:67]
  assign frameBufferDma_clock = clock;
  assign frameBufferDma_reset = reset;
  assign frameBufferDma_io_start = io_enable & io_swap; // @[SpriteFrameBuffer.scala 121:40]
  assign frameBufferDma_io_out_wait_n = ddrArbiter_io_in_1_wait_n; // @[BurstMemIO.scala 156:19 BurstMemArbiter.scala 68:67]
  assign frameBufferDma_io_out_burstDone = ddrArbiter_io_in_1_burstDone; // @[BurstMemIO.scala 156:19 BurstMemArbiter.scala 68:67]
  assign ddrArbiter_clock = clock;
  assign ddrArbiter_reset = reset;
  assign ddrArbiter_io_in_0_rd = lineBufferDma_io_in_rd; // @[BurstMemIO.scala 89:19 90:12]
  assign ddrArbiter_io_in_0_addr = _mem_T_2 + _GEN_2; // @[SpriteFrameBuffer.scala 132:61]
  assign ddrArbiter_io_in_1_wr = frameBufferDma_io_out_wr; // @[BurstMemIO.scala 180:19 181:12]
  assign ddrArbiter_io_in_1_addr = frameBufferDma_io_out_addr + pageFlipper_io_addrWrite; // @[SpriteFrameBuffer.scala 133:37]
  assign ddrArbiter_io_in_1_din = frameBufferDma_io_out_din; // @[BurstMemIO.scala 180:19 187:13]
  assign ddrArbiter_io_in_2_wr = queue_io_out_wr; // @[BurstMemIO.scala 180:19 181:12]
  assign ddrArbiter_io_in_2_addr = queue_io_out_addr + pageFlipper_io_addrWrite; // @[SpriteFrameBuffer.scala 134:28]
  assign ddrArbiter_io_in_2_mask = queue_io_out_mask; // @[BurstMemIO.scala 180:19 186:14]
  assign ddrArbiter_io_in_2_din = queue_io_out_din; // @[BurstMemIO.scala 180:19 187:13]
  assign ddrArbiter_io_out_dout = io_ddr_dout; // @[SpriteFrameBuffer.scala 135:5]
  assign ddrArbiter_io_out_wait_n = io_ddr_wait_n; // @[SpriteFrameBuffer.scala 135:5]
  assign ddrArbiter_io_out_valid = io_ddr_valid; // @[SpriteFrameBuffer.scala 135:5]
  assign ddrArbiter_io_out_burstDone = io_ddr_burstDone; // @[SpriteFrameBuffer.scala 135:5]
  always @(posedge clock) begin
    hBlank_r <= io_video_hBlank; // @[Reg.scala 19:16 20:{18,22}]
    hBlank <= hBlank_r; // @[Reg.scala 19:16 20:{18,22}]
    hBlankRising_REG <= hBlank; // @[Util.scala 158:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hBlank_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  hBlank = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  hBlankRising_REG = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PageFlipper_1(
  input         clock,
  input         reset,
  input         io_mode,
  input         io_swapRead,
  input         io_swapWrite,
  output [31:0] io_addrRead,
  output [31:0] io_addrWrite
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] rdIndexReg; // @[PageFlipper.scala 59:27]
  reg [1:0] wrIndexReg; // @[PageFlipper.scala 60:27]
  wire  _wrIndexReg_T_1 = rdIndexReg == 2'h1; // @[PageFlipper.scala 99:24]
  wire  _wrIndexReg_T_3 = wrIndexReg == 2'h1; // @[PageFlipper.scala 99:39]
  wire  _wrIndexReg_T_6 = wrIndexReg == 2'h0 & rdIndexReg == 2'h1 | wrIndexReg == 2'h1 & rdIndexReg == 2'h0; // @[PageFlipper.scala 99:33]
  wire  _wrIndexReg_T_13 = _wrIndexReg_T_3 & rdIndexReg == 2'h2 | wrIndexReg == 2'h2 & _wrIndexReg_T_1; // @[PageFlipper.scala 100:33]
  wire  _wrIndexReg_T_14 = _wrIndexReg_T_13 ? 1'h0 : 1'h1; // @[Mux.scala 101:16]
  wire [1:0] _wrIndexReg_T_15 = _wrIndexReg_T_6 ? 2'h2 : {{1'd0}, _wrIndexReg_T_14}; // @[Mux.scala 101:16]
  wire  _rdIndexReg_T_6 = rdIndexReg == 2'h0 & wrIndexReg == 2'h1 | rdIndexReg == 2'h1 & wrIndexReg == 2'h0; // @[PageFlipper.scala 99:33]
  wire  _rdIndexReg_T_13 = _wrIndexReg_T_1 & wrIndexReg == 2'h2 | rdIndexReg == 2'h2 & _wrIndexReg_T_3; // @[PageFlipper.scala 100:33]
  wire  _rdIndexReg_T_14 = _rdIndexReg_T_13 ? 1'h0 : 1'h1; // @[Mux.scala 101:16]
  wire [1:0] _rdIndexReg_T_15 = _rdIndexReg_T_6 ? 2'h2 : {{1'd0}, _rdIndexReg_T_14}; // @[Mux.scala 101:16]
  wire [1:0] _GEN_0 = io_swapWrite ? _wrIndexReg_T_15 : wrIndexReg; // @[PageFlipper.scala 68:30 69:18 60:27]
  wire  _wrIndexReg_T_33 = ~wrIndexReg[0]; // @[PageFlipper.scala 75:21]
  wire [12:0] _io_addrRead_T_1 = {11'h120,rdIndexReg}; // @[PageFlipper.scala 80:37]
  wire [12:0] _io_addrWrite_T_1 = {11'h120,wrIndexReg}; // @[PageFlipper.scala 81:38]
  assign io_addrRead = {_io_addrRead_T_1,19'h0}; // @[PageFlipper.scala 80:57]
  assign io_addrWrite = {_io_addrWrite_T_1,19'h0}; // @[PageFlipper.scala 81:58]
  always @(posedge clock) begin
    if (reset) begin // @[PageFlipper.scala 59:27]
      rdIndexReg <= 2'h0; // @[PageFlipper.scala 59:27]
    end else if (io_mode) begin // @[PageFlipper.scala 62:17]
      if (io_swapRead & io_swapWrite) begin // @[PageFlipper.scala 63:39]
        rdIndexReg <= wrIndexReg; // @[PageFlipper.scala 64:18]
      end else if (io_swapRead) begin // @[PageFlipper.scala 66:29]
        rdIndexReg <= _rdIndexReg_T_15; // @[PageFlipper.scala 67:18]
      end
    end else if (io_swapWrite) begin // @[PageFlipper.scala 73:24]
      rdIndexReg <= {{1'd0}, wrIndexReg[0]}; // @[PageFlipper.scala 74:18]
    end
    if (reset) begin // @[PageFlipper.scala 60:27]
      wrIndexReg <= 2'h1; // @[PageFlipper.scala 60:27]
    end else if (io_mode) begin // @[PageFlipper.scala 62:17]
      if (io_swapRead & io_swapWrite) begin // @[PageFlipper.scala 63:39]
        if (_wrIndexReg_T_6) begin // @[Mux.scala 101:16]
          wrIndexReg <= 2'h2;
        end else begin
          wrIndexReg <= {{1'd0}, _wrIndexReg_T_14};
        end
      end else if (!(io_swapRead)) begin // @[PageFlipper.scala 66:29]
        wrIndexReg <= _GEN_0;
      end
    end else if (io_swapWrite) begin // @[PageFlipper.scala 73:24]
      wrIndexReg <= {{1'd0}, _wrIndexReg_T_33}; // @[PageFlipper.scala 75:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rdIndexReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  wrIndexReg = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DualClockFIFO_7(
  input         clock,
  input         io_readClock,
  input         io_deq_ready,
  output        io_deq_valid,
  output [16:0] io_deq_bits_addr,
  output [31:0] io_deq_bits_din,
  output [3:0]  io_deq_bits_mask,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_wr,
  input  [16:0] io_enq_bits_addr,
  input  [31:0] io_enq_bits_din
);
  wire [53:0] fifo_data; // @[DualClockFIFO.scala 74:20]
  wire  fifo_rdclk; // @[DualClockFIFO.scala 74:20]
  wire  fifo_rdreq; // @[DualClockFIFO.scala 74:20]
  wire  fifo_wrclk; // @[DualClockFIFO.scala 74:20]
  wire  fifo_wrreq; // @[DualClockFIFO.scala 74:20]
  wire [53:0] fifo_q; // @[DualClockFIFO.scala 74:20]
  wire  fifo_rdempty; // @[DualClockFIFO.scala 74:20]
  wire  fifo_wrfull; // @[DualClockFIFO.scala 74:20]
  wire [35:0] fifo_io_data_lo = {io_enq_bits_din,4'hf}; // @[DualClockFIFO.scala 80:31]
  wire [17:0] fifo_io_data_hi = {io_enq_bits_wr,io_enq_bits_addr}; // @[DualClockFIFO.scala 80:31]
  wire [53:0] _io_deq_bits_WIRE_1 = fifo_q;
  dual_clock_fifo #(.DATA_WIDTH(54), .DEPTH(16)) fifo ( // @[DualClockFIFO.scala 74:20]
    .data(fifo_data),
    .rdclk(fifo_rdclk),
    .rdreq(fifo_rdreq),
    .wrclk(fifo_wrclk),
    .wrreq(fifo_wrreq),
    .q(fifo_q),
    .rdempty(fifo_rdempty),
    .wrfull(fifo_wrfull)
  );
  assign io_deq_valid = ~fifo_rdempty; // @[DualClockFIFO.scala 85:19]
  assign io_deq_bits_addr = _io_deq_bits_WIRE_1[52:36]; // @[DualClockFIFO.scala 86:36]
  assign io_deq_bits_din = _io_deq_bits_WIRE_1[35:4]; // @[DualClockFIFO.scala 86:36]
  assign io_deq_bits_mask = _io_deq_bits_WIRE_1[3:0]; // @[DualClockFIFO.scala 86:36]
  assign io_enq_ready = ~fifo_wrfull; // @[DualClockFIFO.scala 79:19]
  assign fifo_data = {fifo_io_data_hi,fifo_io_data_lo}; // @[DualClockFIFO.scala 80:31]
  assign fifo_rdclk = io_readClock; // @[DualClockFIFO.scala 83:17]
  assign fifo_rdreq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  assign fifo_wrclk = clock; // @[DualClockFIFO.scala 77:17]
  assign fifo_wrreq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
endmodule
module RequestQueue_1(
  input         clock,
  input         io_enable,
  input         io_readClock,
  input         io_in_wr,
  input  [16:0] io_in_addr,
  input  [31:0] io_in_din,
  output        io_out_wr,
  output [31:0] io_out_addr,
  output [7:0]  io_out_mask,
  output [63:0] io_out_din,
  input         io_out_wait_n
);
  wire  fifo_clock; // @[RequestQueue.scala 70:20]
  wire  fifo_io_readClock; // @[RequestQueue.scala 70:20]
  wire  fifo_io_deq_ready; // @[RequestQueue.scala 70:20]
  wire  fifo_io_deq_valid; // @[RequestQueue.scala 70:20]
  wire [16:0] fifo_io_deq_bits_addr; // @[RequestQueue.scala 70:20]
  wire [31:0] fifo_io_deq_bits_din; // @[RequestQueue.scala 70:20]
  wire [3:0] fifo_io_deq_bits_mask; // @[RequestQueue.scala 70:20]
  wire  fifo_io_enq_ready; // @[RequestQueue.scala 70:20]
  wire  fifo_io_enq_valid; // @[RequestQueue.scala 70:20]
  wire  fifo_io_enq_bits_wr; // @[RequestQueue.scala 70:20]
  wire [16:0] fifo_io_enq_bits_addr; // @[RequestQueue.scala 70:20]
  wire [31:0] fifo_io_enq_bits_din; // @[RequestQueue.scala 70:20]
  wire [18:0] _io_out_addr_T = {fifo_io_deq_bits_addr, 2'h0}; // @[RequestQueue.scala 83:31]
  wire [7:0] _io_out_mask_T_1 = {fifo_io_deq_bits_mask, 4'h0}; // @[RequestQueue.scala 103:54]
  DualClockFIFO_7 fifo ( // @[RequestQueue.scala 70:20]
    .clock(fifo_clock),
    .io_readClock(fifo_io_readClock),
    .io_deq_ready(fifo_io_deq_ready),
    .io_deq_valid(fifo_io_deq_valid),
    .io_deq_bits_addr(fifo_io_deq_bits_addr),
    .io_deq_bits_din(fifo_io_deq_bits_din),
    .io_deq_bits_mask(fifo_io_deq_bits_mask),
    .io_enq_ready(fifo_io_enq_ready),
    .io_enq_valid(fifo_io_enq_valid),
    .io_enq_bits_wr(fifo_io_enq_bits_wr),
    .io_enq_bits_addr(fifo_io_enq_bits_addr),
    .io_enq_bits_din(fifo_io_enq_bits_din)
  );
  assign io_out_wr = io_enable & fifo_io_deq_valid; // @[RequestQueue.scala 79:26]
  assign io_out_addr = {{13'd0}, _io_out_addr_T}; // @[RequestQueue.scala 83:15]
  assign io_out_mask = fifo_io_deq_bits_addr[0] ? _io_out_mask_T_1 : {{4'd0}, fifo_io_deq_bits_mask}; // @[RequestQueue.scala 103:23]
  assign io_out_din = {fifo_io_deq_bits_din,fifo_io_deq_bits_din}; // @[Cat.scala 33:92]
  assign fifo_clock = clock;
  assign fifo_io_readClock = io_readClock; // @[RequestQueue.scala 71:21]
  assign fifo_io_deq_ready = io_out_wait_n; // @[RequestQueue.scala 80:21]
  assign fifo_io_enq_valid = io_in_wr; // @[RequestQueue.scala 74:21]
  assign fifo_io_enq_bits_wr = io_in_wr; // @[WriteRequest.scala 75:19 76:12]
  assign fifo_io_enq_bits_addr = io_in_addr; // @[WriteRequest.scala 75:19 77:14]
  assign fifo_io_enq_bits_din = io_in_din; // @[WriteRequest.scala 75:19 78:13]
endmodule
module SystemFrameBuffer(
  input         clock,
  input         reset,
  input         io_videoClock,
  input         io_enable,
  input         io_rotate,
  input         io_forceBlank,
  input         io_video_vBlank,
  input  [8:0]  io_video_regs_size_x,
  input  [8:0]  io_video_regs_size_y,
  output        io_frameBufferCtrl_enable,
  output [11:0] io_frameBufferCtrl_hSize,
  output [11:0] io_frameBufferCtrl_vSize,
  output [31:0] io_frameBufferCtrl_baseAddr,
  output [13:0] io_frameBufferCtrl_stride,
  input         io_frameBufferCtrl_vBlank,
  input         io_frameBufferCtrl_lowLat,
  output        io_frameBufferCtrl_forceBlank,
  input         io_frameBuffer_wr,
  input  [16:0] io_frameBuffer_addr,
  input  [31:0] io_frameBuffer_din,
  output        io_ddr_wr,
  output [31:0] io_ddr_addr,
  output [7:0]  io_ddr_mask,
  output [63:0] io_ddr_din,
  input         io_ddr_wait_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  pageFlipper_clock; // @[SystemFrameBuffer.scala 80:27]
  wire  pageFlipper_reset; // @[SystemFrameBuffer.scala 80:27]
  wire  pageFlipper_io_mode; // @[SystemFrameBuffer.scala 80:27]
  wire  pageFlipper_io_swapRead; // @[SystemFrameBuffer.scala 80:27]
  wire  pageFlipper_io_swapWrite; // @[SystemFrameBuffer.scala 80:27]
  wire [31:0] pageFlipper_io_addrRead; // @[SystemFrameBuffer.scala 80:27]
  wire [31:0] pageFlipper_io_addrWrite; // @[SystemFrameBuffer.scala 80:27]
  wire  queue_clock; // @[SystemFrameBuffer.scala 98:11]
  wire  queue_io_enable; // @[SystemFrameBuffer.scala 98:11]
  wire  queue_io_readClock; // @[SystemFrameBuffer.scala 98:11]
  wire  queue_io_in_wr; // @[SystemFrameBuffer.scala 98:11]
  wire [16:0] queue_io_in_addr; // @[SystemFrameBuffer.scala 98:11]
  wire [31:0] queue_io_in_din; // @[SystemFrameBuffer.scala 98:11]
  wire  queue_io_out_wr; // @[SystemFrameBuffer.scala 98:11]
  wire [31:0] queue_io_out_addr; // @[SystemFrameBuffer.scala 98:11]
  wire [7:0] queue_io_out_mask; // @[SystemFrameBuffer.scala 98:11]
  wire [63:0] queue_io_out_din; // @[SystemFrameBuffer.scala 98:11]
  wire  queue_io_out_wait_n; // @[SystemFrameBuffer.scala 98:11]
  reg  pageFlipper_io_swapRead_r; // @[Reg.scala 19:16]
  reg  pageFlipper_io_swapRead_r_1; // @[Reg.scala 19:16]
  reg  pageFlipper_io_swapRead_REG; // @[Util.scala 158:44]
  reg  pageFlipper_io_swapWrite_r; // @[Reg.scala 19:16]
  reg  pageFlipper_io_swapWrite_r_1; // @[Reg.scala 19:16]
  reg  pageFlipper_io_swapWrite_REG; // @[Util.scala 158:44]
  wire [8:0] _io_frameBufferCtrl_hSize_T = io_rotate ? io_video_regs_size_y : io_video_regs_size_x; // @[FrameBufferCtrlIO.scala 72:17]
  wire [8:0] _io_frameBufferCtrl_vSize_T = io_rotate ? io_video_regs_size_x : io_video_regs_size_y; // @[FrameBufferCtrlIO.scala 73:17]
  wire [10:0] _io_frameBufferCtrl_stride_T = {io_video_regs_size_y, 2'h0}; // @[FrameBufferCtrlIO.scala 76:34]
  wire [10:0] _io_frameBufferCtrl_stride_T_1 = {io_video_regs_size_x, 2'h0}; // @[FrameBufferCtrlIO.scala 76:46]
  wire [10:0] _io_frameBufferCtrl_stride_T_2 = io_rotate ? _io_frameBufferCtrl_stride_T : _io_frameBufferCtrl_stride_T_1
    ; // @[FrameBufferCtrlIO.scala 76:18]
  PageFlipper_1 pageFlipper ( // @[SystemFrameBuffer.scala 80:27]
    .clock(pageFlipper_clock),
    .reset(pageFlipper_reset),
    .io_mode(pageFlipper_io_mode),
    .io_swapRead(pageFlipper_io_swapRead),
    .io_swapWrite(pageFlipper_io_swapWrite),
    .io_addrRead(pageFlipper_io_addrRead),
    .io_addrWrite(pageFlipper_io_addrWrite)
  );
  RequestQueue_1 queue ( // @[SystemFrameBuffer.scala 98:11]
    .clock(queue_clock),
    .io_enable(queue_io_enable),
    .io_readClock(queue_io_readClock),
    .io_in_wr(queue_io_in_wr),
    .io_in_addr(queue_io_in_addr),
    .io_in_din(queue_io_in_din),
    .io_out_wr(queue_io_out_wr),
    .io_out_addr(queue_io_out_addr),
    .io_out_mask(queue_io_out_mask),
    .io_out_din(queue_io_out_din),
    .io_out_wait_n(queue_io_out_wait_n)
  );
  assign io_frameBufferCtrl_enable = io_enable; // @[FrameBufferCtrlIO.scala 71:17]
  assign io_frameBufferCtrl_hSize = {{3'd0}, _io_frameBufferCtrl_hSize_T}; // @[FrameBufferCtrlIO.scala 72:11]
  assign io_frameBufferCtrl_vSize = {{3'd0}, _io_frameBufferCtrl_vSize_T}; // @[FrameBufferCtrlIO.scala 73:11]
  assign io_frameBufferCtrl_baseAddr = pageFlipper_io_addrRead; // @[FrameBufferCtrlIO.scala 75:19]
  assign io_frameBufferCtrl_stride = {{3'd0}, _io_frameBufferCtrl_stride_T_2}; // @[FrameBufferCtrlIO.scala 76:12]
  assign io_frameBufferCtrl_forceBlank = io_forceBlank; // @[FrameBufferCtrlIO.scala 77:21]
  assign io_ddr_wr = queue_io_out_wr; // @[BurstMemIO.scala 180:19 181:12]
  assign io_ddr_addr = queue_io_out_addr + pageFlipper_io_addrWrite; // @[SystemFrameBuffer.scala 108:26]
  assign io_ddr_mask = queue_io_out_mask; // @[BurstMemIO.scala 180:19 186:14]
  assign io_ddr_din = queue_io_out_din; // @[BurstMemIO.scala 180:19 187:13]
  assign pageFlipper_clock = clock;
  assign pageFlipper_reset = reset;
  assign pageFlipper_io_mode = ~io_frameBufferCtrl_lowLat; // @[SystemFrameBuffer.scala 81:26]
  assign pageFlipper_io_swapRead = pageFlipper_io_swapRead_r_1 & ~pageFlipper_io_swapRead_REG; // @[Util.scala 158:33]
  assign pageFlipper_io_swapWrite = pageFlipper_io_swapWrite_r_1 & ~pageFlipper_io_swapWrite_REG; // @[Util.scala 158:33]
  assign queue_clock = io_videoClock;
  assign queue_io_enable = io_enable; // @[SystemFrameBuffer.scala 106:19]
  assign queue_io_readClock = clock; // @[SystemFrameBuffer.scala 107:22]
  assign queue_io_in_wr = io_frameBuffer_wr; // @[SystemFrameBuffer.scala 111:18]
  assign queue_io_in_addr = io_frameBuffer_addr; // @[SystemFrameBuffer.scala 111:18]
  assign queue_io_in_din = io_frameBuffer_din; // @[SystemFrameBuffer.scala 111:18]
  assign queue_io_out_wait_n = io_ddr_wait_n; // @[BurstMemIO.scala 156:19 SystemFrameBuffer.scala 108:67]
  always @(posedge clock) begin
    pageFlipper_io_swapRead_r <= io_frameBufferCtrl_vBlank; // @[Reg.scala 19:16 20:{18,22}]
    pageFlipper_io_swapRead_r_1 <= pageFlipper_io_swapRead_r; // @[Reg.scala 19:16 20:{18,22}]
    pageFlipper_io_swapRead_REG <= pageFlipper_io_swapRead_r_1; // @[Util.scala 158:44]
    pageFlipper_io_swapWrite_r <= io_video_vBlank; // @[Reg.scala 19:16 20:{18,22}]
    pageFlipper_io_swapWrite_r_1 <= pageFlipper_io_swapWrite_r; // @[Reg.scala 19:16 20:{18,22}]
    pageFlipper_io_swapWrite_REG <= pageFlipper_io_swapWrite_r_1; // @[Util.scala 158:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pageFlipper_io_swapRead_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  pageFlipper_io_swapRead_r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  pageFlipper_io_swapRead_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pageFlipper_io_swapWrite_r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pageFlipper_io_swapWrite_r_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  pageFlipper_io_swapWrite_REG = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cave(
  input         clock,
  input         reset,
  input         cpuClock,
  input         cpuReset,
  input         videoClock,
  input         videoReset,
  input  [3:0]  options_offset_x,
  input  [3:0]  options_offset_y,
  input         options_rotate,
  input         options_compatibility,
  input         options_service,
  input         options_layer_0,
  input         options_layer_1,
  input         options_layer_2,
  input         options_sprite,
  input         options_flip,
  input  [3:0]  options_gameIndex,
  input         player_0_up,
  input         player_0_down,
  input         player_0_left,
  input         player_0_right,
  input  [3:0]  player_0_buttons,
  input         player_0_start,
  input         player_0_coin,
  input         player_0_pause,
  input         player_1_up,
  input         player_1_down,
  input         player_1_left,
  input         player_1_right,
  input  [3:0]  player_1_buttons,
  input         player_1_start,
  input         player_1_coin,
  input         player_1_pause,
  input         ioctl_download,
  input         ioctl_upload,
  input         ioctl_rd,
  input         ioctl_wr,
  output        ioctl_wait_n,
  input  [7:0]  ioctl_index,
  input  [26:0] ioctl_addr,
  output [15:0] ioctl_din,
  input  [15:0] ioctl_dout,
  output        led_power,
  output        led_disk,
  output        led_user,
  output        frameBufferCtrl_enable,
  output [11:0] frameBufferCtrl_hSize,
  output [11:0] frameBufferCtrl_vSize,
  output [4:0]  frameBufferCtrl_format,
  output [31:0] frameBufferCtrl_baseAddr,
  output [13:0] frameBufferCtrl_stride,
  input         frameBufferCtrl_vBlank,
  input         frameBufferCtrl_lowLat,
  output        frameBufferCtrl_forceBlank,
  output        video_clockEnable,
  output        video_displayEnable,
  output [8:0]  video_pos_x,
  output [8:0]  video_pos_y,
  output        video_hSync,
  output        video_vSync,
  output        video_hBlank,
  output        video_vBlank,
  output [8:0]  video_regs_size_x,
  output [8:0]  video_regs_size_y,
  output [8:0]  video_regs_frontPorch_x,
  output [8:0]  video_regs_frontPorch_y,
  output [8:0]  video_regs_retrace_x,
  output [8:0]  video_regs_retrace_y,
  output        video_changeMode,
  output [23:0] rgb,
  output [15:0] audio,
  output        sdram_cke,
  output        sdram_cs_n,
  output        sdram_ras_n,
  output        sdram_cas_n,
  output        sdram_we_n,
  output        sdram_oe_n,
  output [1:0]  sdram_bank,
  output [12:0] sdram_addr,
  output [15:0] sdram_din,
  input  [15:0] sdram_dout,
  output        ddr_rd,
  output        ddr_wr,
  output [31:0] ddr_addr,
  output [7:0]  ddr_mask,
  output [63:0] ddr_din,
  input  [63:0] ddr_dout,
  input         ddr_wait_n,
  input         ddr_valid,
  output [7:0]  ddr_burstLength,
  input         ddr_burstDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  dipsRegs_clock; // @[Cave.scala 112:24]
  wire  dipsRegs_io_mem_wr; // @[Cave.scala 112:24]
  wire [1:0] dipsRegs_io_mem_addr; // @[Cave.scala 112:24]
  wire [15:0] dipsRegs_io_mem_din; // @[Cave.scala 112:24]
  wire [15:0] dipsRegs_io_regs_0; // @[Cave.scala 112:24]
  wire  ddr_1_clock; // @[Cave.scala 118:19]
  wire  ddr_1_reset; // @[Cave.scala 118:19]
  wire  ddr_1_io_mem_rd; // @[Cave.scala 118:19]
  wire  ddr_1_io_mem_wr; // @[Cave.scala 118:19]
  wire [31:0] ddr_1_io_mem_addr; // @[Cave.scala 118:19]
  wire [7:0] ddr_1_io_mem_mask; // @[Cave.scala 118:19]
  wire [63:0] ddr_1_io_mem_din; // @[Cave.scala 118:19]
  wire [63:0] ddr_1_io_mem_dout; // @[Cave.scala 118:19]
  wire  ddr_1_io_mem_wait_n; // @[Cave.scala 118:19]
  wire  ddr_1_io_mem_valid; // @[Cave.scala 118:19]
  wire [7:0] ddr_1_io_mem_burstLength; // @[Cave.scala 118:19]
  wire  ddr_1_io_mem_burstDone; // @[Cave.scala 118:19]
  wire  ddr_1_io_ddr_rd; // @[Cave.scala 118:19]
  wire  ddr_1_io_ddr_wr; // @[Cave.scala 118:19]
  wire [31:0] ddr_1_io_ddr_addr; // @[Cave.scala 118:19]
  wire [7:0] ddr_1_io_ddr_mask; // @[Cave.scala 118:19]
  wire [63:0] ddr_1_io_ddr_din; // @[Cave.scala 118:19]
  wire [63:0] ddr_1_io_ddr_dout; // @[Cave.scala 118:19]
  wire  ddr_1_io_ddr_wait_n; // @[Cave.scala 118:19]
  wire  ddr_1_io_ddr_valid; // @[Cave.scala 118:19]
  wire [7:0] ddr_1_io_ddr_burstLength; // @[Cave.scala 118:19]
  wire  sdram_1_clock; // @[Cave.scala 122:21]
  wire  sdram_1_reset; // @[Cave.scala 122:21]
  wire  sdram_1_io_mem_rd; // @[Cave.scala 122:21]
  wire  sdram_1_io_mem_wr; // @[Cave.scala 122:21]
  wire [24:0] sdram_1_io_mem_addr; // @[Cave.scala 122:21]
  wire [15:0] sdram_1_io_mem_din; // @[Cave.scala 122:21]
  wire [15:0] sdram_1_io_mem_dout; // @[Cave.scala 122:21]
  wire  sdram_1_io_mem_wait_n; // @[Cave.scala 122:21]
  wire  sdram_1_io_mem_valid; // @[Cave.scala 122:21]
  wire  sdram_1_io_mem_burstDone; // @[Cave.scala 122:21]
  wire  sdram_1_io_sdram_cs_n; // @[Cave.scala 122:21]
  wire  sdram_1_io_sdram_ras_n; // @[Cave.scala 122:21]
  wire  sdram_1_io_sdram_cas_n; // @[Cave.scala 122:21]
  wire  sdram_1_io_sdram_we_n; // @[Cave.scala 122:21]
  wire  sdram_1_io_sdram_oe_n; // @[Cave.scala 122:21]
  wire [1:0] sdram_1_io_sdram_bank; // @[Cave.scala 122:21]
  wire [12:0] sdram_1_io_sdram_addr; // @[Cave.scala 122:21]
  wire [15:0] sdram_1_io_sdram_din; // @[Cave.scala 122:21]
  wire [15:0] sdram_1_io_sdram_dout; // @[Cave.scala 122:21]
  wire  memSys_clock; // @[Cave.scala 126:22]
  wire  memSys_reset; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_gameConfig_eepromOffset; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_gameConfig_sound_0_romOffset; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_gameConfig_sound_1_romOffset; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_gameConfig_layer_0_romOffset; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_gameConfig_layer_1_romOffset; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_gameConfig_layer_2_romOffset; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_gameConfig_sprite_romOffset; // @[Cave.scala 126:22]
  wire  memSys_io_prog_rom_wr; // @[Cave.scala 126:22]
  wire [26:0] memSys_io_prog_rom_addr; // @[Cave.scala 126:22]
  wire [15:0] memSys_io_prog_rom_din; // @[Cave.scala 126:22]
  wire  memSys_io_prog_rom_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_prog_nvram_rd; // @[Cave.scala 126:22]
  wire  memSys_io_prog_nvram_wr; // @[Cave.scala 126:22]
  wire [26:0] memSys_io_prog_nvram_addr; // @[Cave.scala 126:22]
  wire [15:0] memSys_io_prog_nvram_din; // @[Cave.scala 126:22]
  wire [15:0] memSys_io_prog_nvram_dout; // @[Cave.scala 126:22]
  wire  memSys_io_prog_nvram_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_prog_nvram_valid; // @[Cave.scala 126:22]
  wire  memSys_io_prog_done; // @[Cave.scala 126:22]
  wire  memSys_io_progRom_rd; // @[Cave.scala 126:22]
  wire [19:0] memSys_io_progRom_addr; // @[Cave.scala 126:22]
  wire [15:0] memSys_io_progRom_dout; // @[Cave.scala 126:22]
  wire  memSys_io_progRom_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_progRom_valid; // @[Cave.scala 126:22]
  wire  memSys_io_eeprom_rd; // @[Cave.scala 126:22]
  wire  memSys_io_eeprom_wr; // @[Cave.scala 126:22]
  wire [6:0] memSys_io_eeprom_addr; // @[Cave.scala 126:22]
  wire [15:0] memSys_io_eeprom_din; // @[Cave.scala 126:22]
  wire [15:0] memSys_io_eeprom_dout; // @[Cave.scala 126:22]
  wire  memSys_io_eeprom_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_eeprom_valid; // @[Cave.scala 126:22]
  wire  memSys_io_soundRom_0_rd; // @[Cave.scala 126:22]
  wire [24:0] memSys_io_soundRom_0_addr; // @[Cave.scala 126:22]
  wire [7:0] memSys_io_soundRom_0_dout; // @[Cave.scala 126:22]
  wire  memSys_io_soundRom_0_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_soundRom_0_valid; // @[Cave.scala 126:22]
  wire  memSys_io_soundRom_1_rd; // @[Cave.scala 126:22]
  wire [24:0] memSys_io_soundRom_1_addr; // @[Cave.scala 126:22]
  wire [7:0] memSys_io_soundRom_1_dout; // @[Cave.scala 126:22]
  wire  memSys_io_soundRom_1_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_soundRom_1_valid; // @[Cave.scala 126:22]
  wire  memSys_io_layerTileRom_0_rd; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_layerTileRom_0_addr; // @[Cave.scala 126:22]
  wire [63:0] memSys_io_layerTileRom_0_dout; // @[Cave.scala 126:22]
  wire  memSys_io_layerTileRom_0_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_layerTileRom_0_valid; // @[Cave.scala 126:22]
  wire  memSys_io_layerTileRom_1_rd; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_layerTileRom_1_addr; // @[Cave.scala 126:22]
  wire [63:0] memSys_io_layerTileRom_1_dout; // @[Cave.scala 126:22]
  wire  memSys_io_layerTileRom_1_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_layerTileRom_1_valid; // @[Cave.scala 126:22]
  wire  memSys_io_layerTileRom_2_rd; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_layerTileRom_2_addr; // @[Cave.scala 126:22]
  wire [63:0] memSys_io_layerTileRom_2_dout; // @[Cave.scala 126:22]
  wire  memSys_io_layerTileRom_2_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_layerTileRom_2_valid; // @[Cave.scala 126:22]
  wire  memSys_io_spriteTileRom_rd; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_spriteTileRom_addr; // @[Cave.scala 126:22]
  wire [63:0] memSys_io_spriteTileRom_dout; // @[Cave.scala 126:22]
  wire  memSys_io_spriteTileRom_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_spriteTileRom_valid; // @[Cave.scala 126:22]
  wire [7:0] memSys_io_spriteTileRom_burstLength; // @[Cave.scala 126:22]
  wire  memSys_io_spriteTileRom_burstDone; // @[Cave.scala 126:22]
  wire  memSys_io_ddr_rd; // @[Cave.scala 126:22]
  wire  memSys_io_ddr_wr; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_ddr_addr; // @[Cave.scala 126:22]
  wire [7:0] memSys_io_ddr_mask; // @[Cave.scala 126:22]
  wire [63:0] memSys_io_ddr_din; // @[Cave.scala 126:22]
  wire [63:0] memSys_io_ddr_dout; // @[Cave.scala 126:22]
  wire  memSys_io_ddr_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_ddr_valid; // @[Cave.scala 126:22]
  wire [7:0] memSys_io_ddr_burstLength; // @[Cave.scala 126:22]
  wire  memSys_io_ddr_burstDone; // @[Cave.scala 126:22]
  wire  memSys_io_sdram_rd; // @[Cave.scala 126:22]
  wire  memSys_io_sdram_wr; // @[Cave.scala 126:22]
  wire [24:0] memSys_io_sdram_addr; // @[Cave.scala 126:22]
  wire [15:0] memSys_io_sdram_din; // @[Cave.scala 126:22]
  wire [15:0] memSys_io_sdram_dout; // @[Cave.scala 126:22]
  wire  memSys_io_sdram_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_sdram_valid; // @[Cave.scala 126:22]
  wire  memSys_io_sdram_burstDone; // @[Cave.scala 126:22]
  wire  memSys_io_spriteFrameBuffer_rd; // @[Cave.scala 126:22]
  wire  memSys_io_spriteFrameBuffer_wr; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_spriteFrameBuffer_addr; // @[Cave.scala 126:22]
  wire [7:0] memSys_io_spriteFrameBuffer_mask; // @[Cave.scala 126:22]
  wire [63:0] memSys_io_spriteFrameBuffer_din; // @[Cave.scala 126:22]
  wire [63:0] memSys_io_spriteFrameBuffer_dout; // @[Cave.scala 126:22]
  wire  memSys_io_spriteFrameBuffer_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_spriteFrameBuffer_valid; // @[Cave.scala 126:22]
  wire [7:0] memSys_io_spriteFrameBuffer_burstLength; // @[Cave.scala 126:22]
  wire  memSys_io_spriteFrameBuffer_burstDone; // @[Cave.scala 126:22]
  wire  memSys_io_systemFrameBuffer_wr; // @[Cave.scala 126:22]
  wire [31:0] memSys_io_systemFrameBuffer_addr; // @[Cave.scala 126:22]
  wire [7:0] memSys_io_systemFrameBuffer_mask; // @[Cave.scala 126:22]
  wire [63:0] memSys_io_systemFrameBuffer_din; // @[Cave.scala 126:22]
  wire  memSys_io_systemFrameBuffer_wait_n; // @[Cave.scala 126:22]
  wire  memSys_io_ready; // @[Cave.scala 126:22]
  wire  videoSys_clock; // @[Cave.scala 135:24]
  wire  videoSys_reset; // @[Cave.scala 135:24]
  wire  videoSys_io_videoClock; // @[Cave.scala 135:24]
  wire  videoSys_io_videoReset; // @[Cave.scala 135:24]
  wire  videoSys_io_prog_video_wr; // @[Cave.scala 135:24]
  wire [26:0] videoSys_io_prog_video_addr; // @[Cave.scala 135:24]
  wire [15:0] videoSys_io_prog_video_din; // @[Cave.scala 135:24]
  wire  videoSys_io_prog_done; // @[Cave.scala 135:24]
  wire [3:0] videoSys_io_options_offset_x; // @[Cave.scala 135:24]
  wire [3:0] videoSys_io_options_offset_y; // @[Cave.scala 135:24]
  wire  videoSys_io_options_compatibility; // @[Cave.scala 135:24]
  wire  videoSys_io_video_clockEnable; // @[Cave.scala 135:24]
  wire  videoSys_io_video_displayEnable; // @[Cave.scala 135:24]
  wire [8:0] videoSys_io_video_pos_x; // @[Cave.scala 135:24]
  wire [8:0] videoSys_io_video_pos_y; // @[Cave.scala 135:24]
  wire  videoSys_io_video_hSync; // @[Cave.scala 135:24]
  wire  videoSys_io_video_vSync; // @[Cave.scala 135:24]
  wire  videoSys_io_video_hBlank; // @[Cave.scala 135:24]
  wire  videoSys_io_video_vBlank; // @[Cave.scala 135:24]
  wire [8:0] videoSys_io_video_regs_size_x; // @[Cave.scala 135:24]
  wire [8:0] videoSys_io_video_regs_size_y; // @[Cave.scala 135:24]
  wire [8:0] videoSys_io_video_regs_frontPorch_x; // @[Cave.scala 135:24]
  wire [8:0] videoSys_io_video_regs_frontPorch_y; // @[Cave.scala 135:24]
  wire [8:0] videoSys_io_video_regs_retrace_x; // @[Cave.scala 135:24]
  wire [8:0] videoSys_io_video_regs_retrace_y; // @[Cave.scala 135:24]
  wire  videoSys_io_video_changeMode; // @[Cave.scala 135:24]
  wire  main_clock; // @[Cave.scala 143:86]
  wire  main_reset; // @[Cave.scala 143:86]
  wire  main_io_videoClock; // @[Cave.scala 143:86]
  wire  main_io_spriteClock; // @[Cave.scala 143:86]
  wire [3:0] main_io_gameIndex; // @[Cave.scala 143:86]
  wire  main_io_options_service; // @[Cave.scala 143:86]
  wire  main_io_player_0_up; // @[Cave.scala 143:86]
  wire  main_io_player_0_down; // @[Cave.scala 143:86]
  wire  main_io_player_0_left; // @[Cave.scala 143:86]
  wire  main_io_player_0_right; // @[Cave.scala 143:86]
  wire [3:0] main_io_player_0_buttons; // @[Cave.scala 143:86]
  wire  main_io_player_0_start; // @[Cave.scala 143:86]
  wire  main_io_player_0_coin; // @[Cave.scala 143:86]
  wire  main_io_player_0_pause; // @[Cave.scala 143:86]
  wire  main_io_player_1_up; // @[Cave.scala 143:86]
  wire  main_io_player_1_down; // @[Cave.scala 143:86]
  wire  main_io_player_1_left; // @[Cave.scala 143:86]
  wire  main_io_player_1_right; // @[Cave.scala 143:86]
  wire [3:0] main_io_player_1_buttons; // @[Cave.scala 143:86]
  wire  main_io_player_1_start; // @[Cave.scala 143:86]
  wire  main_io_player_1_coin; // @[Cave.scala 143:86]
  wire  main_io_player_1_pause; // @[Cave.scala 143:86]
  wire [15:0] main_io_dips_0; // @[Cave.scala 143:86]
  wire  main_io_video_vBlank; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_0_regs_tileSize; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_0_regs_enable; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_0_regs_flipX; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_0_regs_flipY; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_0_regs_rowScrollEnable; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_0_regs_rowSelectEnable; // @[Cave.scala 143:86]
  wire [8:0] main_io_gpuMem_layer_0_regs_scroll_x; // @[Cave.scala 143:86]
  wire [8:0] main_io_gpuMem_layer_0_regs_scroll_y; // @[Cave.scala 143:86]
  wire [11:0] main_io_gpuMem_layer_0_vram8x8_addr; // @[Cave.scala 143:86]
  wire [31:0] main_io_gpuMem_layer_0_vram8x8_dout; // @[Cave.scala 143:86]
  wire [9:0] main_io_gpuMem_layer_0_vram16x16_addr; // @[Cave.scala 143:86]
  wire [31:0] main_io_gpuMem_layer_0_vram16x16_dout; // @[Cave.scala 143:86]
  wire [8:0] main_io_gpuMem_layer_0_lineRam_addr; // @[Cave.scala 143:86]
  wire [31:0] main_io_gpuMem_layer_0_lineRam_dout; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_1_regs_tileSize; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_1_regs_enable; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_1_regs_flipX; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_1_regs_flipY; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_1_regs_rowScrollEnable; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_1_regs_rowSelectEnable; // @[Cave.scala 143:86]
  wire [8:0] main_io_gpuMem_layer_1_regs_scroll_x; // @[Cave.scala 143:86]
  wire [8:0] main_io_gpuMem_layer_1_regs_scroll_y; // @[Cave.scala 143:86]
  wire [11:0] main_io_gpuMem_layer_1_vram8x8_addr; // @[Cave.scala 143:86]
  wire [31:0] main_io_gpuMem_layer_1_vram8x8_dout; // @[Cave.scala 143:86]
  wire [9:0] main_io_gpuMem_layer_1_vram16x16_addr; // @[Cave.scala 143:86]
  wire [31:0] main_io_gpuMem_layer_1_vram16x16_dout; // @[Cave.scala 143:86]
  wire [8:0] main_io_gpuMem_layer_1_lineRam_addr; // @[Cave.scala 143:86]
  wire [31:0] main_io_gpuMem_layer_1_lineRam_dout; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_2_regs_tileSize; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_2_regs_enable; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_2_regs_flipX; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_2_regs_flipY; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_2_regs_rowScrollEnable; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_layer_2_regs_rowSelectEnable; // @[Cave.scala 143:86]
  wire [8:0] main_io_gpuMem_layer_2_regs_scroll_x; // @[Cave.scala 143:86]
  wire [8:0] main_io_gpuMem_layer_2_regs_scroll_y; // @[Cave.scala 143:86]
  wire [11:0] main_io_gpuMem_layer_2_vram8x8_addr; // @[Cave.scala 143:86]
  wire [31:0] main_io_gpuMem_layer_2_vram8x8_dout; // @[Cave.scala 143:86]
  wire [9:0] main_io_gpuMem_layer_2_vram16x16_addr; // @[Cave.scala 143:86]
  wire [31:0] main_io_gpuMem_layer_2_vram16x16_dout; // @[Cave.scala 143:86]
  wire [8:0] main_io_gpuMem_layer_2_lineRam_addr; // @[Cave.scala 143:86]
  wire [31:0] main_io_gpuMem_layer_2_lineRam_dout; // @[Cave.scala 143:86]
  wire [8:0] main_io_gpuMem_sprite_regs_offset_x; // @[Cave.scala 143:86]
  wire [8:0] main_io_gpuMem_sprite_regs_offset_y; // @[Cave.scala 143:86]
  wire [1:0] main_io_gpuMem_sprite_regs_bank; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_sprite_regs_fixed; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_sprite_regs_hFlip; // @[Cave.scala 143:86]
  wire  main_io_gpuMem_sprite_vram_rd; // @[Cave.scala 143:86]
  wire [11:0] main_io_gpuMem_sprite_vram_addr; // @[Cave.scala 143:86]
  wire [127:0] main_io_gpuMem_sprite_vram_dout; // @[Cave.scala 143:86]
  wire [14:0] main_io_gpuMem_paletteRam_addr; // @[Cave.scala 143:86]
  wire [15:0] main_io_gpuMem_paletteRam_dout; // @[Cave.scala 143:86]
  wire  main_io_soundCtrl_oki_0_wr; // @[Cave.scala 143:86]
  wire [15:0] main_io_soundCtrl_oki_0_din; // @[Cave.scala 143:86]
  wire [15:0] main_io_soundCtrl_oki_0_dout; // @[Cave.scala 143:86]
  wire  main_io_soundCtrl_oki_1_wr; // @[Cave.scala 143:86]
  wire [15:0] main_io_soundCtrl_oki_1_din; // @[Cave.scala 143:86]
  wire [15:0] main_io_soundCtrl_oki_1_dout; // @[Cave.scala 143:86]
  wire  main_io_soundCtrl_nmk_wr; // @[Cave.scala 143:86]
  wire [22:0] main_io_soundCtrl_nmk_addr; // @[Cave.scala 143:86]
  wire [15:0] main_io_soundCtrl_nmk_din; // @[Cave.scala 143:86]
  wire  main_io_soundCtrl_ymz_rd; // @[Cave.scala 143:86]
  wire  main_io_soundCtrl_ymz_wr; // @[Cave.scala 143:86]
  wire [22:0] main_io_soundCtrl_ymz_addr; // @[Cave.scala 143:86]
  wire [15:0] main_io_soundCtrl_ymz_din; // @[Cave.scala 143:86]
  wire [15:0] main_io_soundCtrl_ymz_dout; // @[Cave.scala 143:86]
  wire  main_io_soundCtrl_req; // @[Cave.scala 143:86]
  wire [15:0] main_io_soundCtrl_data; // @[Cave.scala 143:86]
  wire  main_io_soundCtrl_irq; // @[Cave.scala 143:86]
  wire  main_io_progRom_rd; // @[Cave.scala 143:86]
  wire [19:0] main_io_progRom_addr; // @[Cave.scala 143:86]
  wire [15:0] main_io_progRom_dout; // @[Cave.scala 143:86]
  wire  main_io_progRom_valid; // @[Cave.scala 143:86]
  wire  main_io_eeprom_rd; // @[Cave.scala 143:86]
  wire  main_io_eeprom_wr; // @[Cave.scala 143:86]
  wire [6:0] main_io_eeprom_addr; // @[Cave.scala 143:86]
  wire [15:0] main_io_eeprom_din; // @[Cave.scala 143:86]
  wire [15:0] main_io_eeprom_dout; // @[Cave.scala 143:86]
  wire  main_io_eeprom_wait_n; // @[Cave.scala 143:86]
  wire  main_io_eeprom_valid; // @[Cave.scala 143:86]
  wire  main_io_spriteFrameBufferSwap; // @[Cave.scala 143:86]
  wire  main_io_progRom_freezer_clock; // @[Crossing.scala 213:25]
  wire  main_io_progRom_freezer_reset; // @[Crossing.scala 213:25]
  wire  main_io_progRom_freezer_io_targetClock; // @[Crossing.scala 213:25]
  wire  main_io_progRom_freezer_io_in_rd; // @[Crossing.scala 213:25]
  wire [19:0] main_io_progRom_freezer_io_in_addr; // @[Crossing.scala 213:25]
  wire [15:0] main_io_progRom_freezer_io_in_dout; // @[Crossing.scala 213:25]
  wire  main_io_progRom_freezer_io_in_valid; // @[Crossing.scala 213:25]
  wire  main_io_progRom_freezer_io_out_rd; // @[Crossing.scala 213:25]
  wire [19:0] main_io_progRom_freezer_io_out_addr; // @[Crossing.scala 213:25]
  wire [15:0] main_io_progRom_freezer_io_out_dout; // @[Crossing.scala 213:25]
  wire  main_io_progRom_freezer_io_out_wait_n; // @[Crossing.scala 213:25]
  wire  main_io_progRom_freezer_io_out_valid; // @[Crossing.scala 213:25]
  wire  main_io_eeprom_freezer_clock; // @[Crossing.scala 226:25]
  wire  main_io_eeprom_freezer_reset; // @[Crossing.scala 226:25]
  wire  main_io_eeprom_freezer_io_targetClock; // @[Crossing.scala 226:25]
  wire  main_io_eeprom_freezer_io_in_rd; // @[Crossing.scala 226:25]
  wire  main_io_eeprom_freezer_io_in_wr; // @[Crossing.scala 226:25]
  wire [6:0] main_io_eeprom_freezer_io_in_addr; // @[Crossing.scala 226:25]
  wire [15:0] main_io_eeprom_freezer_io_in_din; // @[Crossing.scala 226:25]
  wire [15:0] main_io_eeprom_freezer_io_in_dout; // @[Crossing.scala 226:25]
  wire  main_io_eeprom_freezer_io_in_wait_n; // @[Crossing.scala 226:25]
  wire  main_io_eeprom_freezer_io_in_valid; // @[Crossing.scala 226:25]
  wire  main_io_eeprom_freezer_io_out_rd; // @[Crossing.scala 226:25]
  wire  main_io_eeprom_freezer_io_out_wr; // @[Crossing.scala 226:25]
  wire [6:0] main_io_eeprom_freezer_io_out_addr; // @[Crossing.scala 226:25]
  wire [15:0] main_io_eeprom_freezer_io_out_din; // @[Crossing.scala 226:25]
  wire [15:0] main_io_eeprom_freezer_io_out_dout; // @[Crossing.scala 226:25]
  wire  main_io_eeprom_freezer_io_out_wait_n; // @[Crossing.scala 226:25]
  wire  main_io_eeprom_freezer_io_out_valid; // @[Crossing.scala 226:25]
  wire  sound_clock; // @[Cave.scala 155:87]
  wire  sound_reset; // @[Cave.scala 155:87]
  wire  sound_io_ctrl_oki_0_wr; // @[Cave.scala 155:87]
  wire [15:0] sound_io_ctrl_oki_0_din; // @[Cave.scala 155:87]
  wire [15:0] sound_io_ctrl_oki_0_dout; // @[Cave.scala 155:87]
  wire  sound_io_ctrl_oki_1_wr; // @[Cave.scala 155:87]
  wire [15:0] sound_io_ctrl_oki_1_din; // @[Cave.scala 155:87]
  wire [15:0] sound_io_ctrl_oki_1_dout; // @[Cave.scala 155:87]
  wire  sound_io_ctrl_nmk_wr; // @[Cave.scala 155:87]
  wire [22:0] sound_io_ctrl_nmk_addr; // @[Cave.scala 155:87]
  wire [15:0] sound_io_ctrl_nmk_din; // @[Cave.scala 155:87]
  wire  sound_io_ctrl_ymz_rd; // @[Cave.scala 155:87]
  wire  sound_io_ctrl_ymz_wr; // @[Cave.scala 155:87]
  wire [22:0] sound_io_ctrl_ymz_addr; // @[Cave.scala 155:87]
  wire [15:0] sound_io_ctrl_ymz_din; // @[Cave.scala 155:87]
  wire [15:0] sound_io_ctrl_ymz_dout; // @[Cave.scala 155:87]
  wire  sound_io_ctrl_req; // @[Cave.scala 155:87]
  wire [15:0] sound_io_ctrl_data; // @[Cave.scala 155:87]
  wire  sound_io_ctrl_irq; // @[Cave.scala 155:87]
  wire [3:0] sound_io_gameIndex; // @[Cave.scala 155:87]
  wire [1:0] sound_io_gameConfig_sound_0_device; // @[Cave.scala 155:87]
  wire  sound_io_rom_0_rd; // @[Cave.scala 155:87]
  wire [24:0] sound_io_rom_0_addr; // @[Cave.scala 155:87]
  wire [7:0] sound_io_rom_0_dout; // @[Cave.scala 155:87]
  wire  sound_io_rom_0_wait_n; // @[Cave.scala 155:87]
  wire  sound_io_rom_0_valid; // @[Cave.scala 155:87]
  wire [24:0] sound_io_rom_1_addr; // @[Cave.scala 155:87]
  wire [7:0] sound_io_rom_1_dout; // @[Cave.scala 155:87]
  wire  sound_io_rom_1_valid; // @[Cave.scala 155:87]
  wire [15:0] sound_io_audio; // @[Cave.scala 155:87]
  wire  sound_io_rom_0_freezer_clock; // @[Crossing.scala 213:25]
  wire  sound_io_rom_0_freezer_reset; // @[Crossing.scala 213:25]
  wire  sound_io_rom_0_freezer_io_targetClock; // @[Crossing.scala 213:25]
  wire  sound_io_rom_0_freezer_io_in_rd; // @[Crossing.scala 213:25]
  wire [24:0] sound_io_rom_0_freezer_io_in_addr; // @[Crossing.scala 213:25]
  wire [7:0] sound_io_rom_0_freezer_io_in_dout; // @[Crossing.scala 213:25]
  wire  sound_io_rom_0_freezer_io_in_wait_n; // @[Crossing.scala 213:25]
  wire  sound_io_rom_0_freezer_io_in_valid; // @[Crossing.scala 213:25]
  wire  sound_io_rom_0_freezer_io_out_rd; // @[Crossing.scala 213:25]
  wire [24:0] sound_io_rom_0_freezer_io_out_addr; // @[Crossing.scala 213:25]
  wire [7:0] sound_io_rom_0_freezer_io_out_dout; // @[Crossing.scala 213:25]
  wire  sound_io_rom_0_freezer_io_out_wait_n; // @[Crossing.scala 213:25]
  wire  sound_io_rom_0_freezer_io_out_valid; // @[Crossing.scala 213:25]
  wire  sound_io_rom_1_freezer_clock; // @[Crossing.scala 213:25]
  wire  sound_io_rom_1_freezer_reset; // @[Crossing.scala 213:25]
  wire  sound_io_rom_1_freezer_io_targetClock; // @[Crossing.scala 213:25]
  wire  sound_io_rom_1_freezer_io_in_rd; // @[Crossing.scala 213:25]
  wire [24:0] sound_io_rom_1_freezer_io_in_addr; // @[Crossing.scala 213:25]
  wire [7:0] sound_io_rom_1_freezer_io_in_dout; // @[Crossing.scala 213:25]
  wire  sound_io_rom_1_freezer_io_in_wait_n; // @[Crossing.scala 213:25]
  wire  sound_io_rom_1_freezer_io_in_valid; // @[Crossing.scala 213:25]
  wire  sound_io_rom_1_freezer_io_out_rd; // @[Crossing.scala 213:25]
  wire [24:0] sound_io_rom_1_freezer_io_out_addr; // @[Crossing.scala 213:25]
  wire [7:0] sound_io_rom_1_freezer_io_out_dout; // @[Crossing.scala 213:25]
  wire  sound_io_rom_1_freezer_io_out_wait_n; // @[Crossing.scala 213:25]
  wire  sound_io_rom_1_freezer_io_out_valid; // @[Crossing.scala 213:25]
  wire  gpu_clock; // @[Cave.scala 163:19]
  wire  gpu_reset; // @[Cave.scala 163:19]
  wire  gpu_io_videoClock; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_0_enable; // @[Cave.scala 163:19]
  wire [1:0] gpu_io_layerCtrl_0_format; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_0_regs_tileSize; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_0_regs_enable; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_0_regs_flipX; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_0_regs_flipY; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_0_regs_rowScrollEnable; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_0_regs_rowSelectEnable; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_layerCtrl_0_regs_scroll_x; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_layerCtrl_0_regs_scroll_y; // @[Cave.scala 163:19]
  wire [11:0] gpu_io_layerCtrl_0_vram8x8_addr; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_layerCtrl_0_vram8x8_dout; // @[Cave.scala 163:19]
  wire [9:0] gpu_io_layerCtrl_0_vram16x16_addr; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_layerCtrl_0_vram16x16_dout; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_layerCtrl_0_lineRam_addr; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_layerCtrl_0_lineRam_dout; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_0_tileRom_rd; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_layerCtrl_0_tileRom_addr; // @[Cave.scala 163:19]
  wire [63:0] gpu_io_layerCtrl_0_tileRom_dout; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_1_enable; // @[Cave.scala 163:19]
  wire [1:0] gpu_io_layerCtrl_1_format; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_1_regs_tileSize; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_1_regs_enable; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_1_regs_flipX; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_1_regs_flipY; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_1_regs_rowScrollEnable; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_1_regs_rowSelectEnable; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_layerCtrl_1_regs_scroll_x; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_layerCtrl_1_regs_scroll_y; // @[Cave.scala 163:19]
  wire [11:0] gpu_io_layerCtrl_1_vram8x8_addr; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_layerCtrl_1_vram8x8_dout; // @[Cave.scala 163:19]
  wire [9:0] gpu_io_layerCtrl_1_vram16x16_addr; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_layerCtrl_1_vram16x16_dout; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_layerCtrl_1_lineRam_addr; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_layerCtrl_1_lineRam_dout; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_1_tileRom_rd; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_layerCtrl_1_tileRom_addr; // @[Cave.scala 163:19]
  wire [63:0] gpu_io_layerCtrl_1_tileRom_dout; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_2_enable; // @[Cave.scala 163:19]
  wire [1:0] gpu_io_layerCtrl_2_format; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_2_regs_tileSize; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_2_regs_enable; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_2_regs_flipX; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_2_regs_flipY; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_2_regs_rowScrollEnable; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_2_regs_rowSelectEnable; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_layerCtrl_2_regs_scroll_x; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_layerCtrl_2_regs_scroll_y; // @[Cave.scala 163:19]
  wire [11:0] gpu_io_layerCtrl_2_vram8x8_addr; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_layerCtrl_2_vram8x8_dout; // @[Cave.scala 163:19]
  wire [9:0] gpu_io_layerCtrl_2_vram16x16_addr; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_layerCtrl_2_vram16x16_dout; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_layerCtrl_2_lineRam_addr; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_layerCtrl_2_lineRam_dout; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_2_tileRom_rd; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_layerCtrl_2_tileRom_addr; // @[Cave.scala 163:19]
  wire [63:0] gpu_io_layerCtrl_2_tileRom_dout; // @[Cave.scala 163:19]
  wire  gpu_io_spriteCtrl_enable; // @[Cave.scala 163:19]
  wire [1:0] gpu_io_spriteCtrl_format; // @[Cave.scala 163:19]
  wire  gpu_io_spriteCtrl_start; // @[Cave.scala 163:19]
  wire  gpu_io_spriteCtrl_zoom; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_spriteCtrl_regs_offset_x; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_spriteCtrl_regs_offset_y; // @[Cave.scala 163:19]
  wire [1:0] gpu_io_spriteCtrl_regs_bank; // @[Cave.scala 163:19]
  wire  gpu_io_spriteCtrl_regs_fixed; // @[Cave.scala 163:19]
  wire  gpu_io_spriteCtrl_regs_hFlip; // @[Cave.scala 163:19]
  wire  gpu_io_spriteCtrl_vram_rd; // @[Cave.scala 163:19]
  wire [11:0] gpu_io_spriteCtrl_vram_addr; // @[Cave.scala 163:19]
  wire [127:0] gpu_io_spriteCtrl_vram_dout; // @[Cave.scala 163:19]
  wire  gpu_io_spriteCtrl_tileRom_rd; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_spriteCtrl_tileRom_addr; // @[Cave.scala 163:19]
  wire [63:0] gpu_io_spriteCtrl_tileRom_dout; // @[Cave.scala 163:19]
  wire  gpu_io_spriteCtrl_tileRom_wait_n; // @[Cave.scala 163:19]
  wire  gpu_io_spriteCtrl_tileRom_valid; // @[Cave.scala 163:19]
  wire [7:0] gpu_io_spriteCtrl_tileRom_burstLength; // @[Cave.scala 163:19]
  wire  gpu_io_spriteCtrl_tileRom_burstDone; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_gameConfig_granularity; // @[Cave.scala 163:19]
  wire [1:0] gpu_io_gameConfig_layer_0_paletteBank; // @[Cave.scala 163:19]
  wire [1:0] gpu_io_gameConfig_layer_1_paletteBank; // @[Cave.scala 163:19]
  wire [1:0] gpu_io_gameConfig_layer_2_paletteBank; // @[Cave.scala 163:19]
  wire  gpu_io_options_rotate; // @[Cave.scala 163:19]
  wire  gpu_io_options_flip; // @[Cave.scala 163:19]
  wire  gpu_io_video_clockEnable; // @[Cave.scala 163:19]
  wire  gpu_io_video_displayEnable; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_video_pos_x; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_video_pos_y; // @[Cave.scala 163:19]
  wire  gpu_io_video_vBlank; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_video_regs_size_x; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_video_regs_size_y; // @[Cave.scala 163:19]
  wire [8:0] gpu_io_spriteLineBuffer_addr; // @[Cave.scala 163:19]
  wire [15:0] gpu_io_spriteLineBuffer_dout; // @[Cave.scala 163:19]
  wire  gpu_io_spriteFrameBuffer_wr; // @[Cave.scala 163:19]
  wire [16:0] gpu_io_spriteFrameBuffer_addr; // @[Cave.scala 163:19]
  wire [15:0] gpu_io_spriteFrameBuffer_din; // @[Cave.scala 163:19]
  wire  gpu_io_spriteFrameBuffer_wait_n; // @[Cave.scala 163:19]
  wire  gpu_io_systemFrameBuffer_wr; // @[Cave.scala 163:19]
  wire [16:0] gpu_io_systemFrameBuffer_addr; // @[Cave.scala 163:19]
  wire [31:0] gpu_io_systemFrameBuffer_din; // @[Cave.scala 163:19]
  wire [14:0] gpu_io_paletteRam_addr; // @[Cave.scala 163:19]
  wire [15:0] gpu_io_paletteRam_dout; // @[Cave.scala 163:19]
  wire [23:0] gpu_io_rgb; // @[Cave.scala 163:19]
  wire  gpu_io_layerCtrl_0_tileRom_crossing_clock; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_0_tileRom_crossing_io_targetClock; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_0_tileRom_crossing_io_in_rd; // @[Crossing.scala 200:26]
  wire [31:0] gpu_io_layerCtrl_0_tileRom_crossing_io_in_addr; // @[Crossing.scala 200:26]
  wire [63:0] gpu_io_layerCtrl_0_tileRom_crossing_io_in_dout; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_0_tileRom_crossing_io_out_rd; // @[Crossing.scala 200:26]
  wire [31:0] gpu_io_layerCtrl_0_tileRom_crossing_io_out_addr; // @[Crossing.scala 200:26]
  wire [63:0] gpu_io_layerCtrl_0_tileRom_crossing_io_out_dout; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_0_tileRom_crossing_io_out_wait_n; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_0_tileRom_crossing_io_out_valid; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_1_tileRom_crossing_clock; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_1_tileRom_crossing_io_targetClock; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_1_tileRom_crossing_io_in_rd; // @[Crossing.scala 200:26]
  wire [31:0] gpu_io_layerCtrl_1_tileRom_crossing_io_in_addr; // @[Crossing.scala 200:26]
  wire [63:0] gpu_io_layerCtrl_1_tileRom_crossing_io_in_dout; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_1_tileRom_crossing_io_out_rd; // @[Crossing.scala 200:26]
  wire [31:0] gpu_io_layerCtrl_1_tileRom_crossing_io_out_addr; // @[Crossing.scala 200:26]
  wire [63:0] gpu_io_layerCtrl_1_tileRom_crossing_io_out_dout; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_1_tileRom_crossing_io_out_wait_n; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_1_tileRom_crossing_io_out_valid; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_2_tileRom_crossing_clock; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_2_tileRom_crossing_io_targetClock; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_2_tileRom_crossing_io_in_rd; // @[Crossing.scala 200:26]
  wire [31:0] gpu_io_layerCtrl_2_tileRom_crossing_io_in_addr; // @[Crossing.scala 200:26]
  wire [63:0] gpu_io_layerCtrl_2_tileRom_crossing_io_in_dout; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_2_tileRom_crossing_io_out_rd; // @[Crossing.scala 200:26]
  wire [31:0] gpu_io_layerCtrl_2_tileRom_crossing_io_out_addr; // @[Crossing.scala 200:26]
  wire [63:0] gpu_io_layerCtrl_2_tileRom_crossing_io_out_dout; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_2_tileRom_crossing_io_out_wait_n; // @[Crossing.scala 200:26]
  wire  gpu_io_layerCtrl_2_tileRom_crossing_io_out_valid; // @[Crossing.scala 200:26]
  wire  spriteFrameBuffer_clock; // @[Cave.scala 187:33]
  wire  spriteFrameBuffer_reset; // @[Cave.scala 187:33]
  wire  spriteFrameBuffer_io_videoClock; // @[Cave.scala 187:33]
  wire  spriteFrameBuffer_io_enable; // @[Cave.scala 187:33]
  wire  spriteFrameBuffer_io_swap; // @[Cave.scala 187:33]
  wire [8:0] spriteFrameBuffer_io_video_pos_y; // @[Cave.scala 187:33]
  wire  spriteFrameBuffer_io_video_hBlank; // @[Cave.scala 187:33]
  wire [8:0] spriteFrameBuffer_io_lineBuffer_addr; // @[Cave.scala 187:33]
  wire [15:0] spriteFrameBuffer_io_lineBuffer_dout; // @[Cave.scala 187:33]
  wire  spriteFrameBuffer_io_frameBuffer_wr; // @[Cave.scala 187:33]
  wire [16:0] spriteFrameBuffer_io_frameBuffer_addr; // @[Cave.scala 187:33]
  wire [15:0] spriteFrameBuffer_io_frameBuffer_din; // @[Cave.scala 187:33]
  wire  spriteFrameBuffer_io_frameBuffer_wait_n; // @[Cave.scala 187:33]
  wire  spriteFrameBuffer_io_ddr_rd; // @[Cave.scala 187:33]
  wire  spriteFrameBuffer_io_ddr_wr; // @[Cave.scala 187:33]
  wire [31:0] spriteFrameBuffer_io_ddr_addr; // @[Cave.scala 187:33]
  wire [7:0] spriteFrameBuffer_io_ddr_mask; // @[Cave.scala 187:33]
  wire [63:0] spriteFrameBuffer_io_ddr_din; // @[Cave.scala 187:33]
  wire [63:0] spriteFrameBuffer_io_ddr_dout; // @[Cave.scala 187:33]
  wire  spriteFrameBuffer_io_ddr_wait_n; // @[Cave.scala 187:33]
  wire  spriteFrameBuffer_io_ddr_valid; // @[Cave.scala 187:33]
  wire [7:0] spriteFrameBuffer_io_ddr_burstLength; // @[Cave.scala 187:33]
  wire  spriteFrameBuffer_io_ddr_burstDone; // @[Cave.scala 187:33]
  wire  systemFrameBuffer_clock; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_reset; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_io_videoClock; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_io_enable; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_io_rotate; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_io_forceBlank; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_io_video_vBlank; // @[Cave.scala 197:33]
  wire [8:0] systemFrameBuffer_io_video_regs_size_x; // @[Cave.scala 197:33]
  wire [8:0] systemFrameBuffer_io_video_regs_size_y; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_io_frameBufferCtrl_enable; // @[Cave.scala 197:33]
  wire [11:0] systemFrameBuffer_io_frameBufferCtrl_hSize; // @[Cave.scala 197:33]
  wire [11:0] systemFrameBuffer_io_frameBufferCtrl_vSize; // @[Cave.scala 197:33]
  wire [31:0] systemFrameBuffer_io_frameBufferCtrl_baseAddr; // @[Cave.scala 197:33]
  wire [13:0] systemFrameBuffer_io_frameBufferCtrl_stride; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_io_frameBufferCtrl_vBlank; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_io_frameBufferCtrl_lowLat; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_io_frameBufferCtrl_forceBlank; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_io_frameBuffer_wr; // @[Cave.scala 197:33]
  wire [16:0] systemFrameBuffer_io_frameBuffer_addr; // @[Cave.scala 197:33]
  wire [31:0] systemFrameBuffer_io_frameBuffer_din; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_io_ddr_wr; // @[Cave.scala 197:33]
  wire [31:0] systemFrameBuffer_io_ddr_addr; // @[Cave.scala 197:33]
  wire [7:0] systemFrameBuffer_io_ddr_mask; // @[Cave.scala 197:33]
  wire [63:0] systemFrameBuffer_io_ddr_din; // @[Cave.scala 197:33]
  wire  systemFrameBuffer_io_ddr_wait_n; // @[Cave.scala 197:33]
  reg  vBlank_r; // @[Reg.scala 19:16]
  reg  vBlank; // @[Reg.scala 19:16]
  reg  vBlankFalling_REG; // @[Util.scala 165:45]
  reg [3:0] gameIndexReg; // @[Cave.scala 95:18]
  reg  gameIndexReg_latched; // @[Cave.scala 96:26]
  wire  _GEN_3 = ioctl_download & ioctl_wr & ioctl_index == 8'h1 | gameIndexReg_latched; // @[Cave.scala 97:85 99:15 96:26]
  reg  gameIndexReg_REG; // @[Util.scala 165:45]
  wire  _gameIndexReg_T_4 = ~ioctl_download & gameIndexReg_REG; // @[Util.scala 165:35]
  wire  _GEN_5 = _gameIndexReg_T_4 & ~gameIndexReg_latched | _GEN_3; // @[Cave.scala 101:55 103:15]
  wire [8:0] _gameConfig_T_1_granularity = 4'h1 == gameIndexReg ? 9'h100 : 9'h10; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_1_layer_2_format = 4'h1 == gameIndexReg ? 2'h3 : 2'h0; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_1_layer_2_romOffset = 4'h1 == gameIndexReg ? 32'h900080 : 32'h0; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_1_layer_2_paletteBank = 4'h1 == gameIndexReg ? 2'h1 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_1_sprite_format = 4'h1 == gameIndexReg ? 2'h2 : 2'h1; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_1_sprite_romOffset = 4'h1 == gameIndexReg ? 32'hb00080 : 32'h900080; // @[Mux.scala 81:58]
  wire  _gameConfig_T_1_sprite_zoom = 4'h1 == gameIndexReg ? 1'h0 : 1'h1; // @[Mux.scala 81:58]
  wire [8:0] _gameConfig_T_3_granularity = 4'h2 == gameIndexReg ? 9'h10 : _gameConfig_T_1_granularity; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_3_eepromOffset = 4'h2 == gameIndexReg ? 32'h80000 : 32'h100000; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_3_sound_0_device = 4'h2 == gameIndexReg ? 2'h2 : 2'h1; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_3_sound_0_romOffset = 4'h2 == gameIndexReg ? 32'h80080 : 32'h100080; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_3_sound_1_romOffset = 4'h2 == gameIndexReg ? 32'h280080 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_3_layer_0_romOffset = 4'h2 == gameIndexReg ? 32'h380080 : 32'h500080; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_3_layer_1_romOffset = 4'h2 == gameIndexReg ? 32'h480080 : 32'h700080; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_3_layer_2_format = 4'h2 == gameIndexReg ? 2'h1 : _gameConfig_T_1_layer_2_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_3_layer_2_romOffset = 4'h2 == gameIndexReg ? 32'h580080 : _gameConfig_T_1_layer_2_romOffset; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_3_layer_2_paletteBank = 4'h2 == gameIndexReg ? 2'h1 : _gameConfig_T_1_layer_2_paletteBank; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_3_sprite_format = 4'h2 == gameIndexReg ? 2'h2 : _gameConfig_T_1_sprite_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_3_sprite_romOffset = 4'h2 == gameIndexReg ? 32'h5c0080 : _gameConfig_T_1_sprite_romOffset; // @[Mux.scala 81:58]
  wire  _gameConfig_T_3_sprite_zoom = 4'h2 == gameIndexReg ? 1'h0 : _gameConfig_T_1_sprite_zoom; // @[Mux.scala 81:58]
  wire [8:0] _gameConfig_T_5_granularity = 4'h3 == gameIndexReg ? 9'h100 : _gameConfig_T_3_granularity; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_5_eepromOffset = 4'h3 == gameIndexReg ? 32'h100000 : _gameConfig_T_3_eepromOffset; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_5_sound_0_device = 4'h3 == gameIndexReg ? 2'h1 : _gameConfig_T_3_sound_0_device; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_5_sound_0_romOffset = 4'h3 == gameIndexReg ? 32'h100080 : _gameConfig_T_3_sound_0_romOffset; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_5_sound_1_romOffset = 4'h3 == gameIndexReg ? 32'h0 : _gameConfig_T_3_sound_1_romOffset; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_5_layer_0_format = 4'h3 == gameIndexReg ? 2'h3 : 2'h1; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_5_layer_0_romOffset = 4'h3 == gameIndexReg ? 32'h500080 : _gameConfig_T_3_layer_0_romOffset; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_5_layer_1_romOffset = 4'h3 == gameIndexReg ? 32'hd00080 : _gameConfig_T_3_layer_1_romOffset; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_5_layer_2_format = 4'h3 == gameIndexReg ? 2'h3 : _gameConfig_T_3_layer_2_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_5_layer_2_romOffset = 4'h3 == gameIndexReg ? 32'h1500080 : _gameConfig_T_3_layer_2_romOffset
    ; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_5_layer_2_paletteBank = 4'h3 == gameIndexReg ? 2'h1 : _gameConfig_T_3_layer_2_paletteBank; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_5_sprite_format = 4'h3 == gameIndexReg ? 2'h3 : _gameConfig_T_3_sprite_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_5_sprite_romOffset = 4'h3 == gameIndexReg ? 32'h1900080 : _gameConfig_T_3_sprite_romOffset; // @[Mux.scala 81:58]
  wire [8:0] _gameConfig_T_7_granularity = 4'h6 == gameIndexReg ? 9'h100 : _gameConfig_T_5_granularity; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_7_eepromOffset = 4'h6 == gameIndexReg ? 32'h0 : _gameConfig_T_5_eepromOffset; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_7_sound_0_device = 4'h6 == gameIndexReg ? 2'h1 : _gameConfig_T_5_sound_0_device; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_7_sound_0_romOffset = 4'h6 == gameIndexReg ? 32'h100000 : _gameConfig_T_5_sound_0_romOffset; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_7_sound_1_romOffset = 4'h6 == gameIndexReg ? 32'h0 : _gameConfig_T_5_sound_1_romOffset; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_7_layer_0_format = 4'h6 == gameIndexReg ? 2'h3 : _gameConfig_T_5_layer_0_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_7_layer_0_romOffset = 4'h6 == gameIndexReg ? 32'hd00000 : _gameConfig_T_5_layer_0_romOffset; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_7_layer_1_romOffset = 4'h6 == gameIndexReg ? 32'h1100000 : _gameConfig_T_5_layer_1_romOffset
    ; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_7_layer_2_format = 4'h6 == gameIndexReg ? 2'h3 : _gameConfig_T_5_layer_2_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_7_layer_2_romOffset = 4'h6 == gameIndexReg ? 32'h1500000 : _gameConfig_T_5_layer_2_romOffset
    ; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_7_layer_2_paletteBank = 4'h6 == gameIndexReg ? 2'h1 : _gameConfig_T_5_layer_2_paletteBank; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_7_sprite_format = 4'h6 == gameIndexReg ? 2'h1 : _gameConfig_T_5_sprite_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_7_sprite_romOffset = 4'h6 == gameIndexReg ? 32'h1900000 : _gameConfig_T_5_sprite_romOffset; // @[Mux.scala 81:58]
  wire [8:0] _gameConfig_T_9_granularity = 4'h5 == gameIndexReg ? 9'h100 : _gameConfig_T_7_granularity; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_9_eepromOffset = 4'h5 == gameIndexReg ? 32'h100000 : _gameConfig_T_7_eepromOffset; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_9_sound_0_device = 4'h5 == gameIndexReg ? 2'h1 : _gameConfig_T_7_sound_0_device; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_9_sound_0_romOffset = 4'h5 == gameIndexReg ? 32'h100080 : _gameConfig_T_7_sound_0_romOffset; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_9_sound_1_romOffset = 4'h5 == gameIndexReg ? 32'h0 : _gameConfig_T_7_sound_1_romOffset; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_9_layer_0_format = 4'h5 == gameIndexReg ? 2'h3 : _gameConfig_T_7_layer_0_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_9_layer_0_romOffset = 4'h5 == gameIndexReg ? 32'h500080 : _gameConfig_T_7_layer_0_romOffset; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_9_layer_1_romOffset = 4'h5 == gameIndexReg ? 32'hd00080 : _gameConfig_T_7_layer_1_romOffset; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_9_layer_2_format = 4'h5 == gameIndexReg ? 2'h3 : _gameConfig_T_7_layer_2_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_9_layer_2_romOffset = 4'h5 == gameIndexReg ? 32'h1100080 : _gameConfig_T_7_layer_2_romOffset
    ; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_9_layer_2_paletteBank = 4'h5 == gameIndexReg ? 2'h1 : _gameConfig_T_7_layer_2_paletteBank; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_9_sprite_format = 4'h5 == gameIndexReg ? 2'h3 : _gameConfig_T_7_sprite_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_9_sprite_romOffset = 4'h5 == gameIndexReg ? 32'h1500080 : _gameConfig_T_7_sprite_romOffset; // @[Mux.scala 81:58]
  wire [8:0] _gameConfig_T_11_granularity = 4'h7 == gameIndexReg ? 9'h10 : _gameConfig_T_9_granularity; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_11_eepromOffset = 4'h7 == gameIndexReg ? 32'h100000 : _gameConfig_T_9_eepromOffset; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_11_sound_0_device = 4'h7 == gameIndexReg ? 2'h3 : _gameConfig_T_9_sound_0_device; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_11_sound_0_romOffset = 4'h7 == gameIndexReg ? 32'h100080 : _gameConfig_T_9_sound_0_romOffset
    ; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_11_sound_1_romOffset = 4'h7 == gameIndexReg ? 32'h140080 : _gameConfig_T_9_sound_1_romOffset
    ; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_11_layer_0_format = 4'h7 == gameIndexReg ? 2'h1 : _gameConfig_T_9_layer_0_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_11_layer_0_romOffset = 4'h7 == gameIndexReg ? 32'h1c0080 : _gameConfig_T_9_layer_0_romOffset
    ; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_11_layer_0_paletteBank = 4'h7 == gameIndexReg ? 2'h0 : 2'h1; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_11_layer_1_romOffset = 4'h7 == gameIndexReg ? 32'h240080 : _gameConfig_T_9_layer_1_romOffset
    ; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_11_layer_2_format = 4'h7 == gameIndexReg ? 2'h1 : _gameConfig_T_9_layer_2_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_11_layer_2_romOffset = 4'h7 == gameIndexReg ? 32'h2c0080 : _gameConfig_T_9_layer_2_romOffset
    ; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_11_layer_2_paletteBank = 4'h7 == gameIndexReg ? 2'h0 : _gameConfig_T_9_layer_2_paletteBank; // @[Mux.scala 81:58]
  wire [1:0] _gameConfig_T_11_sprite_format = 4'h7 == gameIndexReg ? 2'h1 : _gameConfig_T_9_sprite_format; // @[Mux.scala 81:58]
  wire [31:0] _gameConfig_T_11_sprite_romOffset = 4'h7 == gameIndexReg ? 32'h340080 : _gameConfig_T_9_sprite_romOffset; // @[Mux.scala 81:58]
  wire  dipsRegs_io_mem_writeEnable = ioctl_download & ioctl_index == 8'hfe & ~(|ioctl_addr[26:3]); // @[IOCTL.scala 94:68]
  wire  _memSys_io_prog_rom_writeEnable_T = ioctl_index == 8'h0; // @[IOCTL.scala 67:46]
  wire  memSys_io_prog_rom_writeEnable = ioctl_download & ioctl_index == 8'h0; // @[IOCTL.scala 67:32]
  wire  memSys_io_prog_rom_mem_wait_n = memSys_io_prog_rom_wait_n; // @[IOCTL.scala 68:19 Cave.scala 128:22]
  wire  _GEN_7 = memSys_io_prog_rom_writeEnable ? memSys_io_prog_rom_mem_wait_n : 1'h1; // @[IOCTL.scala 70:{23,32}]
  wire  _memSys_io_prog_nvram_readEnable_T = ioctl_index == 8'h2; // @[IOCTL.scala 79:43]
  wire  memSys_io_prog_nvram_readEnable = ioctl_upload & ioctl_index == 8'h2; // @[IOCTL.scala 79:29]
  wire  memSys_io_prog_nvram_writeEnable = ioctl_download & _memSys_io_prog_nvram_readEnable_T; // @[IOCTL.scala 80:32]
  wire  memSys_io_prog_nvram_mem_wait_n = memSys_io_prog_nvram_wait_n; // @[IOCTL.scala 81:19 Cave.scala 129:24]
  wire  _GEN_8 = memSys_io_prog_nvram_readEnable | memSys_io_prog_nvram_writeEnable ? memSys_io_prog_nvram_mem_wait_n :
    _GEN_7; // @[IOCTL.scala 84:{37,46}]
  reg [15:0] memSys_io_prog_nvram_view__ioctl_din_r; // @[Reg.scala 19:16]
  wire  memSys_io_prog_nvram_mem_valid = memSys_io_prog_nvram_valid; // @[IOCTL.scala 81:19 Cave.scala 129:24]
  wire [15:0] memSys_io_prog_nvram_mem_dout = memSys_io_prog_nvram_dout; // @[IOCTL.scala 81:19 Cave.scala 129:24]
  reg  memSys_io_prog_done_REG; // @[Util.scala 165:45]
  wire  _memSys_io_prog_done_T_1 = ~ioctl_download & memSys_io_prog_done_REG; // @[Util.scala 165:35]
  wire  _videoSys_io_prog_video_writeEnable_T = ioctl_index == 8'h3; // @[IOCTL.scala 106:46]
  wire  videoSys_io_prog_video_writeEnable = ioctl_download & ioctl_index == 8'h3; // @[IOCTL.scala 106:32]
  reg  videoSys_io_prog_done_REG; // @[Util.scala 165:45]
  wire  _videoSys_io_prog_done_T_1 = ~ioctl_download & videoSys_io_prog_done_REG; // @[Util.scala 165:35]
  wire  _T = ~memSys_io_ready; // @[Cave.scala 143:60]
  RegisterFile dipsRegs ( // @[Cave.scala 112:24]
    .clock(dipsRegs_clock),
    .io_mem_wr(dipsRegs_io_mem_wr),
    .io_mem_addr(dipsRegs_io_mem_addr),
    .io_mem_din(dipsRegs_io_mem_din),
    .io_regs_0(dipsRegs_io_regs_0)
  );
  DDR ddr_1 ( // @[Cave.scala 118:19]
    .clock(ddr_1_clock),
    .reset(ddr_1_reset),
    .io_mem_rd(ddr_1_io_mem_rd),
    .io_mem_wr(ddr_1_io_mem_wr),
    .io_mem_addr(ddr_1_io_mem_addr),
    .io_mem_mask(ddr_1_io_mem_mask),
    .io_mem_din(ddr_1_io_mem_din),
    .io_mem_dout(ddr_1_io_mem_dout),
    .io_mem_wait_n(ddr_1_io_mem_wait_n),
    .io_mem_valid(ddr_1_io_mem_valid),
    .io_mem_burstLength(ddr_1_io_mem_burstLength),
    .io_mem_burstDone(ddr_1_io_mem_burstDone),
    .io_ddr_rd(ddr_1_io_ddr_rd),
    .io_ddr_wr(ddr_1_io_ddr_wr),
    .io_ddr_addr(ddr_1_io_ddr_addr),
    .io_ddr_mask(ddr_1_io_ddr_mask),
    .io_ddr_din(ddr_1_io_ddr_din),
    .io_ddr_dout(ddr_1_io_ddr_dout),
    .io_ddr_wait_n(ddr_1_io_ddr_wait_n),
    .io_ddr_valid(ddr_1_io_ddr_valid),
    .io_ddr_burstLength(ddr_1_io_ddr_burstLength)
  );
  SDRAM sdram_1 ( // @[Cave.scala 122:21]
    .clock(sdram_1_clock),
    .reset(sdram_1_reset),
    .io_mem_rd(sdram_1_io_mem_rd),
    .io_mem_wr(sdram_1_io_mem_wr),
    .io_mem_addr(sdram_1_io_mem_addr),
    .io_mem_din(sdram_1_io_mem_din),
    .io_mem_dout(sdram_1_io_mem_dout),
    .io_mem_wait_n(sdram_1_io_mem_wait_n),
    .io_mem_valid(sdram_1_io_mem_valid),
    .io_mem_burstDone(sdram_1_io_mem_burstDone),
    .io_sdram_cs_n(sdram_1_io_sdram_cs_n),
    .io_sdram_ras_n(sdram_1_io_sdram_ras_n),
    .io_sdram_cas_n(sdram_1_io_sdram_cas_n),
    .io_sdram_we_n(sdram_1_io_sdram_we_n),
    .io_sdram_oe_n(sdram_1_io_sdram_oe_n),
    .io_sdram_bank(sdram_1_io_sdram_bank),
    .io_sdram_addr(sdram_1_io_sdram_addr),
    .io_sdram_din(sdram_1_io_sdram_din),
    .io_sdram_dout(sdram_1_io_sdram_dout)
  );
  MemSys memSys ( // @[Cave.scala 126:22]
    .clock(memSys_clock),
    .reset(memSys_reset),
    .io_gameConfig_eepromOffset(memSys_io_gameConfig_eepromOffset),
    .io_gameConfig_sound_0_romOffset(memSys_io_gameConfig_sound_0_romOffset),
    .io_gameConfig_sound_1_romOffset(memSys_io_gameConfig_sound_1_romOffset),
    .io_gameConfig_layer_0_romOffset(memSys_io_gameConfig_layer_0_romOffset),
    .io_gameConfig_layer_1_romOffset(memSys_io_gameConfig_layer_1_romOffset),
    .io_gameConfig_layer_2_romOffset(memSys_io_gameConfig_layer_2_romOffset),
    .io_gameConfig_sprite_romOffset(memSys_io_gameConfig_sprite_romOffset),
    .io_prog_rom_wr(memSys_io_prog_rom_wr),
    .io_prog_rom_addr(memSys_io_prog_rom_addr),
    .io_prog_rom_din(memSys_io_prog_rom_din),
    .io_prog_rom_wait_n(memSys_io_prog_rom_wait_n),
    .io_prog_nvram_rd(memSys_io_prog_nvram_rd),
    .io_prog_nvram_wr(memSys_io_prog_nvram_wr),
    .io_prog_nvram_addr(memSys_io_prog_nvram_addr),
    .io_prog_nvram_din(memSys_io_prog_nvram_din),
    .io_prog_nvram_dout(memSys_io_prog_nvram_dout),
    .io_prog_nvram_wait_n(memSys_io_prog_nvram_wait_n),
    .io_prog_nvram_valid(memSys_io_prog_nvram_valid),
    .io_prog_done(memSys_io_prog_done),
    .io_progRom_rd(memSys_io_progRom_rd),
    .io_progRom_addr(memSys_io_progRom_addr),
    .io_progRom_dout(memSys_io_progRom_dout),
    .io_progRom_wait_n(memSys_io_progRom_wait_n),
    .io_progRom_valid(memSys_io_progRom_valid),
    .io_eeprom_rd(memSys_io_eeprom_rd),
    .io_eeprom_wr(memSys_io_eeprom_wr),
    .io_eeprom_addr(memSys_io_eeprom_addr),
    .io_eeprom_din(memSys_io_eeprom_din),
    .io_eeprom_dout(memSys_io_eeprom_dout),
    .io_eeprom_wait_n(memSys_io_eeprom_wait_n),
    .io_eeprom_valid(memSys_io_eeprom_valid),
    .io_soundRom_0_rd(memSys_io_soundRom_0_rd),
    .io_soundRom_0_addr(memSys_io_soundRom_0_addr),
    .io_soundRom_0_dout(memSys_io_soundRom_0_dout),
    .io_soundRom_0_wait_n(memSys_io_soundRom_0_wait_n),
    .io_soundRom_0_valid(memSys_io_soundRom_0_valid),
    .io_soundRom_1_rd(memSys_io_soundRom_1_rd),
    .io_soundRom_1_addr(memSys_io_soundRom_1_addr),
    .io_soundRom_1_dout(memSys_io_soundRom_1_dout),
    .io_soundRom_1_wait_n(memSys_io_soundRom_1_wait_n),
    .io_soundRom_1_valid(memSys_io_soundRom_1_valid),
    .io_layerTileRom_0_rd(memSys_io_layerTileRom_0_rd),
    .io_layerTileRom_0_addr(memSys_io_layerTileRom_0_addr),
    .io_layerTileRom_0_dout(memSys_io_layerTileRom_0_dout),
    .io_layerTileRom_0_wait_n(memSys_io_layerTileRom_0_wait_n),
    .io_layerTileRom_0_valid(memSys_io_layerTileRom_0_valid),
    .io_layerTileRom_1_rd(memSys_io_layerTileRom_1_rd),
    .io_layerTileRom_1_addr(memSys_io_layerTileRom_1_addr),
    .io_layerTileRom_1_dout(memSys_io_layerTileRom_1_dout),
    .io_layerTileRom_1_wait_n(memSys_io_layerTileRom_1_wait_n),
    .io_layerTileRom_1_valid(memSys_io_layerTileRom_1_valid),
    .io_layerTileRom_2_rd(memSys_io_layerTileRom_2_rd),
    .io_layerTileRom_2_addr(memSys_io_layerTileRom_2_addr),
    .io_layerTileRom_2_dout(memSys_io_layerTileRom_2_dout),
    .io_layerTileRom_2_wait_n(memSys_io_layerTileRom_2_wait_n),
    .io_layerTileRom_2_valid(memSys_io_layerTileRom_2_valid),
    .io_spriteTileRom_rd(memSys_io_spriteTileRom_rd),
    .io_spriteTileRom_addr(memSys_io_spriteTileRom_addr),
    .io_spriteTileRom_dout(memSys_io_spriteTileRom_dout),
    .io_spriteTileRom_wait_n(memSys_io_spriteTileRom_wait_n),
    .io_spriteTileRom_valid(memSys_io_spriteTileRom_valid),
    .io_spriteTileRom_burstLength(memSys_io_spriteTileRom_burstLength),
    .io_spriteTileRom_burstDone(memSys_io_spriteTileRom_burstDone),
    .io_ddr_rd(memSys_io_ddr_rd),
    .io_ddr_wr(memSys_io_ddr_wr),
    .io_ddr_addr(memSys_io_ddr_addr),
    .io_ddr_mask(memSys_io_ddr_mask),
    .io_ddr_din(memSys_io_ddr_din),
    .io_ddr_dout(memSys_io_ddr_dout),
    .io_ddr_wait_n(memSys_io_ddr_wait_n),
    .io_ddr_valid(memSys_io_ddr_valid),
    .io_ddr_burstLength(memSys_io_ddr_burstLength),
    .io_ddr_burstDone(memSys_io_ddr_burstDone),
    .io_sdram_rd(memSys_io_sdram_rd),
    .io_sdram_wr(memSys_io_sdram_wr),
    .io_sdram_addr(memSys_io_sdram_addr),
    .io_sdram_din(memSys_io_sdram_din),
    .io_sdram_dout(memSys_io_sdram_dout),
    .io_sdram_wait_n(memSys_io_sdram_wait_n),
    .io_sdram_valid(memSys_io_sdram_valid),
    .io_sdram_burstDone(memSys_io_sdram_burstDone),
    .io_spriteFrameBuffer_rd(memSys_io_spriteFrameBuffer_rd),
    .io_spriteFrameBuffer_wr(memSys_io_spriteFrameBuffer_wr),
    .io_spriteFrameBuffer_addr(memSys_io_spriteFrameBuffer_addr),
    .io_spriteFrameBuffer_mask(memSys_io_spriteFrameBuffer_mask),
    .io_spriteFrameBuffer_din(memSys_io_spriteFrameBuffer_din),
    .io_spriteFrameBuffer_dout(memSys_io_spriteFrameBuffer_dout),
    .io_spriteFrameBuffer_wait_n(memSys_io_spriteFrameBuffer_wait_n),
    .io_spriteFrameBuffer_valid(memSys_io_spriteFrameBuffer_valid),
    .io_spriteFrameBuffer_burstLength(memSys_io_spriteFrameBuffer_burstLength),
    .io_spriteFrameBuffer_burstDone(memSys_io_spriteFrameBuffer_burstDone),
    .io_systemFrameBuffer_wr(memSys_io_systemFrameBuffer_wr),
    .io_systemFrameBuffer_addr(memSys_io_systemFrameBuffer_addr),
    .io_systemFrameBuffer_mask(memSys_io_systemFrameBuffer_mask),
    .io_systemFrameBuffer_din(memSys_io_systemFrameBuffer_din),
    .io_systemFrameBuffer_wait_n(memSys_io_systemFrameBuffer_wait_n),
    .io_ready(memSys_io_ready)
  );
  VideoSys videoSys ( // @[Cave.scala 135:24]
    .clock(videoSys_clock),
    .reset(videoSys_reset),
    .io_videoClock(videoSys_io_videoClock),
    .io_videoReset(videoSys_io_videoReset),
    .io_prog_video_wr(videoSys_io_prog_video_wr),
    .io_prog_video_addr(videoSys_io_prog_video_addr),
    .io_prog_video_din(videoSys_io_prog_video_din),
    .io_prog_done(videoSys_io_prog_done),
    .io_options_offset_x(videoSys_io_options_offset_x),
    .io_options_offset_y(videoSys_io_options_offset_y),
    .io_options_compatibility(videoSys_io_options_compatibility),
    .io_video_clockEnable(videoSys_io_video_clockEnable),
    .io_video_displayEnable(videoSys_io_video_displayEnable),
    .io_video_pos_x(videoSys_io_video_pos_x),
    .io_video_pos_y(videoSys_io_video_pos_y),
    .io_video_hSync(videoSys_io_video_hSync),
    .io_video_vSync(videoSys_io_video_vSync),
    .io_video_hBlank(videoSys_io_video_hBlank),
    .io_video_vBlank(videoSys_io_video_vBlank),
    .io_video_regs_size_x(videoSys_io_video_regs_size_x),
    .io_video_regs_size_y(videoSys_io_video_regs_size_y),
    .io_video_regs_frontPorch_x(videoSys_io_video_regs_frontPorch_x),
    .io_video_regs_frontPorch_y(videoSys_io_video_regs_frontPorch_y),
    .io_video_regs_retrace_x(videoSys_io_video_regs_retrace_x),
    .io_video_regs_retrace_y(videoSys_io_video_regs_retrace_y),
    .io_video_changeMode(videoSys_io_video_changeMode)
  );
  Main main ( // @[Cave.scala 143:86]
    .clock(main_clock),
    .reset(main_reset),
    .io_videoClock(main_io_videoClock),
    .io_spriteClock(main_io_spriteClock),
    .io_gameIndex(main_io_gameIndex),
    .io_options_service(main_io_options_service),
    .io_player_0_up(main_io_player_0_up),
    .io_player_0_down(main_io_player_0_down),
    .io_player_0_left(main_io_player_0_left),
    .io_player_0_right(main_io_player_0_right),
    .io_player_0_buttons(main_io_player_0_buttons),
    .io_player_0_start(main_io_player_0_start),
    .io_player_0_coin(main_io_player_0_coin),
    .io_player_0_pause(main_io_player_0_pause),
    .io_player_1_up(main_io_player_1_up),
    .io_player_1_down(main_io_player_1_down),
    .io_player_1_left(main_io_player_1_left),
    .io_player_1_right(main_io_player_1_right),
    .io_player_1_buttons(main_io_player_1_buttons),
    .io_player_1_start(main_io_player_1_start),
    .io_player_1_coin(main_io_player_1_coin),
    .io_player_1_pause(main_io_player_1_pause),
    .io_dips_0(main_io_dips_0),
    .io_video_vBlank(main_io_video_vBlank),
    .io_gpuMem_layer_0_regs_tileSize(main_io_gpuMem_layer_0_regs_tileSize),
    .io_gpuMem_layer_0_regs_enable(main_io_gpuMem_layer_0_regs_enable),
    .io_gpuMem_layer_0_regs_flipX(main_io_gpuMem_layer_0_regs_flipX),
    .io_gpuMem_layer_0_regs_flipY(main_io_gpuMem_layer_0_regs_flipY),
    .io_gpuMem_layer_0_regs_rowScrollEnable(main_io_gpuMem_layer_0_regs_rowScrollEnable),
    .io_gpuMem_layer_0_regs_rowSelectEnable(main_io_gpuMem_layer_0_regs_rowSelectEnable),
    .io_gpuMem_layer_0_regs_scroll_x(main_io_gpuMem_layer_0_regs_scroll_x),
    .io_gpuMem_layer_0_regs_scroll_y(main_io_gpuMem_layer_0_regs_scroll_y),
    .io_gpuMem_layer_0_vram8x8_addr(main_io_gpuMem_layer_0_vram8x8_addr),
    .io_gpuMem_layer_0_vram8x8_dout(main_io_gpuMem_layer_0_vram8x8_dout),
    .io_gpuMem_layer_0_vram16x16_addr(main_io_gpuMem_layer_0_vram16x16_addr),
    .io_gpuMem_layer_0_vram16x16_dout(main_io_gpuMem_layer_0_vram16x16_dout),
    .io_gpuMem_layer_0_lineRam_addr(main_io_gpuMem_layer_0_lineRam_addr),
    .io_gpuMem_layer_0_lineRam_dout(main_io_gpuMem_layer_0_lineRam_dout),
    .io_gpuMem_layer_1_regs_tileSize(main_io_gpuMem_layer_1_regs_tileSize),
    .io_gpuMem_layer_1_regs_enable(main_io_gpuMem_layer_1_regs_enable),
    .io_gpuMem_layer_1_regs_flipX(main_io_gpuMem_layer_1_regs_flipX),
    .io_gpuMem_layer_1_regs_flipY(main_io_gpuMem_layer_1_regs_flipY),
    .io_gpuMem_layer_1_regs_rowScrollEnable(main_io_gpuMem_layer_1_regs_rowScrollEnable),
    .io_gpuMem_layer_1_regs_rowSelectEnable(main_io_gpuMem_layer_1_regs_rowSelectEnable),
    .io_gpuMem_layer_1_regs_scroll_x(main_io_gpuMem_layer_1_regs_scroll_x),
    .io_gpuMem_layer_1_regs_scroll_y(main_io_gpuMem_layer_1_regs_scroll_y),
    .io_gpuMem_layer_1_vram8x8_addr(main_io_gpuMem_layer_1_vram8x8_addr),
    .io_gpuMem_layer_1_vram8x8_dout(main_io_gpuMem_layer_1_vram8x8_dout),
    .io_gpuMem_layer_1_vram16x16_addr(main_io_gpuMem_layer_1_vram16x16_addr),
    .io_gpuMem_layer_1_vram16x16_dout(main_io_gpuMem_layer_1_vram16x16_dout),
    .io_gpuMem_layer_1_lineRam_addr(main_io_gpuMem_layer_1_lineRam_addr),
    .io_gpuMem_layer_1_lineRam_dout(main_io_gpuMem_layer_1_lineRam_dout),
    .io_gpuMem_layer_2_regs_tileSize(main_io_gpuMem_layer_2_regs_tileSize),
    .io_gpuMem_layer_2_regs_enable(main_io_gpuMem_layer_2_regs_enable),
    .io_gpuMem_layer_2_regs_flipX(main_io_gpuMem_layer_2_regs_flipX),
    .io_gpuMem_layer_2_regs_flipY(main_io_gpuMem_layer_2_regs_flipY),
    .io_gpuMem_layer_2_regs_rowScrollEnable(main_io_gpuMem_layer_2_regs_rowScrollEnable),
    .io_gpuMem_layer_2_regs_rowSelectEnable(main_io_gpuMem_layer_2_regs_rowSelectEnable),
    .io_gpuMem_layer_2_regs_scroll_x(main_io_gpuMem_layer_2_regs_scroll_x),
    .io_gpuMem_layer_2_regs_scroll_y(main_io_gpuMem_layer_2_regs_scroll_y),
    .io_gpuMem_layer_2_vram8x8_addr(main_io_gpuMem_layer_2_vram8x8_addr),
    .io_gpuMem_layer_2_vram8x8_dout(main_io_gpuMem_layer_2_vram8x8_dout),
    .io_gpuMem_layer_2_vram16x16_addr(main_io_gpuMem_layer_2_vram16x16_addr),
    .io_gpuMem_layer_2_vram16x16_dout(main_io_gpuMem_layer_2_vram16x16_dout),
    .io_gpuMem_layer_2_lineRam_addr(main_io_gpuMem_layer_2_lineRam_addr),
    .io_gpuMem_layer_2_lineRam_dout(main_io_gpuMem_layer_2_lineRam_dout),
    .io_gpuMem_sprite_regs_offset_x(main_io_gpuMem_sprite_regs_offset_x),
    .io_gpuMem_sprite_regs_offset_y(main_io_gpuMem_sprite_regs_offset_y),
    .io_gpuMem_sprite_regs_bank(main_io_gpuMem_sprite_regs_bank),
    .io_gpuMem_sprite_regs_fixed(main_io_gpuMem_sprite_regs_fixed),
    .io_gpuMem_sprite_regs_hFlip(main_io_gpuMem_sprite_regs_hFlip),
    .io_gpuMem_sprite_vram_rd(main_io_gpuMem_sprite_vram_rd),
    .io_gpuMem_sprite_vram_addr(main_io_gpuMem_sprite_vram_addr),
    .io_gpuMem_sprite_vram_dout(main_io_gpuMem_sprite_vram_dout),
    .io_gpuMem_paletteRam_addr(main_io_gpuMem_paletteRam_addr),
    .io_gpuMem_paletteRam_dout(main_io_gpuMem_paletteRam_dout),
    .io_soundCtrl_oki_0_wr(main_io_soundCtrl_oki_0_wr),
    .io_soundCtrl_oki_0_din(main_io_soundCtrl_oki_0_din),
    .io_soundCtrl_oki_0_dout(main_io_soundCtrl_oki_0_dout),
    .io_soundCtrl_oki_1_wr(main_io_soundCtrl_oki_1_wr),
    .io_soundCtrl_oki_1_din(main_io_soundCtrl_oki_1_din),
    .io_soundCtrl_oki_1_dout(main_io_soundCtrl_oki_1_dout),
    .io_soundCtrl_nmk_wr(main_io_soundCtrl_nmk_wr),
    .io_soundCtrl_nmk_addr(main_io_soundCtrl_nmk_addr),
    .io_soundCtrl_nmk_din(main_io_soundCtrl_nmk_din),
    .io_soundCtrl_ymz_rd(main_io_soundCtrl_ymz_rd),
    .io_soundCtrl_ymz_wr(main_io_soundCtrl_ymz_wr),
    .io_soundCtrl_ymz_addr(main_io_soundCtrl_ymz_addr),
    .io_soundCtrl_ymz_din(main_io_soundCtrl_ymz_din),
    .io_soundCtrl_ymz_dout(main_io_soundCtrl_ymz_dout),
    .io_soundCtrl_req(main_io_soundCtrl_req),
    .io_soundCtrl_data(main_io_soundCtrl_data),
    .io_soundCtrl_irq(main_io_soundCtrl_irq),
    .io_progRom_rd(main_io_progRom_rd),
    .io_progRom_addr(main_io_progRom_addr),
    .io_progRom_dout(main_io_progRom_dout),
    .io_progRom_valid(main_io_progRom_valid),
    .io_eeprom_rd(main_io_eeprom_rd),
    .io_eeprom_wr(main_io_eeprom_wr),
    .io_eeprom_addr(main_io_eeprom_addr),
    .io_eeprom_din(main_io_eeprom_din),
    .io_eeprom_dout(main_io_eeprom_dout),
    .io_eeprom_wait_n(main_io_eeprom_wait_n),
    .io_eeprom_valid(main_io_eeprom_valid),
    .io_spriteFrameBufferSwap(main_io_spriteFrameBufferSwap)
  );
  ReadDataFreezer main_io_progRom_freezer ( // @[Crossing.scala 213:25]
    .clock(main_io_progRom_freezer_clock),
    .reset(main_io_progRom_freezer_reset),
    .io_targetClock(main_io_progRom_freezer_io_targetClock),
    .io_in_rd(main_io_progRom_freezer_io_in_rd),
    .io_in_addr(main_io_progRom_freezer_io_in_addr),
    .io_in_dout(main_io_progRom_freezer_io_in_dout),
    .io_in_valid(main_io_progRom_freezer_io_in_valid),
    .io_out_rd(main_io_progRom_freezer_io_out_rd),
    .io_out_addr(main_io_progRom_freezer_io_out_addr),
    .io_out_dout(main_io_progRom_freezer_io_out_dout),
    .io_out_wait_n(main_io_progRom_freezer_io_out_wait_n),
    .io_out_valid(main_io_progRom_freezer_io_out_valid)
  );
  DataFreezer main_io_eeprom_freezer ( // @[Crossing.scala 226:25]
    .clock(main_io_eeprom_freezer_clock),
    .reset(main_io_eeprom_freezer_reset),
    .io_targetClock(main_io_eeprom_freezer_io_targetClock),
    .io_in_rd(main_io_eeprom_freezer_io_in_rd),
    .io_in_wr(main_io_eeprom_freezer_io_in_wr),
    .io_in_addr(main_io_eeprom_freezer_io_in_addr),
    .io_in_din(main_io_eeprom_freezer_io_in_din),
    .io_in_dout(main_io_eeprom_freezer_io_in_dout),
    .io_in_wait_n(main_io_eeprom_freezer_io_in_wait_n),
    .io_in_valid(main_io_eeprom_freezer_io_in_valid),
    .io_out_rd(main_io_eeprom_freezer_io_out_rd),
    .io_out_wr(main_io_eeprom_freezer_io_out_wr),
    .io_out_addr(main_io_eeprom_freezer_io_out_addr),
    .io_out_din(main_io_eeprom_freezer_io_out_din),
    .io_out_dout(main_io_eeprom_freezer_io_out_dout),
    .io_out_wait_n(main_io_eeprom_freezer_io_out_wait_n),
    .io_out_valid(main_io_eeprom_freezer_io_out_valid)
  );
  Sound sound ( // @[Cave.scala 155:87]
    .clock(sound_clock),
    .reset(sound_reset),
    .io_ctrl_oki_0_wr(sound_io_ctrl_oki_0_wr),
    .io_ctrl_oki_0_din(sound_io_ctrl_oki_0_din),
    .io_ctrl_oki_0_dout(sound_io_ctrl_oki_0_dout),
    .io_ctrl_oki_1_wr(sound_io_ctrl_oki_1_wr),
    .io_ctrl_oki_1_din(sound_io_ctrl_oki_1_din),
    .io_ctrl_oki_1_dout(sound_io_ctrl_oki_1_dout),
    .io_ctrl_nmk_wr(sound_io_ctrl_nmk_wr),
    .io_ctrl_nmk_addr(sound_io_ctrl_nmk_addr),
    .io_ctrl_nmk_din(sound_io_ctrl_nmk_din),
    .io_ctrl_ymz_rd(sound_io_ctrl_ymz_rd),
    .io_ctrl_ymz_wr(sound_io_ctrl_ymz_wr),
    .io_ctrl_ymz_addr(sound_io_ctrl_ymz_addr),
    .io_ctrl_ymz_din(sound_io_ctrl_ymz_din),
    .io_ctrl_ymz_dout(sound_io_ctrl_ymz_dout),
    .io_ctrl_req(sound_io_ctrl_req),
    .io_ctrl_data(sound_io_ctrl_data),
    .io_ctrl_irq(sound_io_ctrl_irq),
    .io_gameIndex(sound_io_gameIndex),
    .io_gameConfig_sound_0_device(sound_io_gameConfig_sound_0_device),
    .io_rom_0_rd(sound_io_rom_0_rd),
    .io_rom_0_addr(sound_io_rom_0_addr),
    .io_rom_0_dout(sound_io_rom_0_dout),
    .io_rom_0_wait_n(sound_io_rom_0_wait_n),
    .io_rom_0_valid(sound_io_rom_0_valid),
    .io_rom_1_addr(sound_io_rom_1_addr),
    .io_rom_1_dout(sound_io_rom_1_dout),
    .io_rom_1_valid(sound_io_rom_1_valid),
    .io_audio(sound_io_audio)
  );
  ReadDataFreezer_1 sound_io_rom_0_freezer ( // @[Crossing.scala 213:25]
    .clock(sound_io_rom_0_freezer_clock),
    .reset(sound_io_rom_0_freezer_reset),
    .io_targetClock(sound_io_rom_0_freezer_io_targetClock),
    .io_in_rd(sound_io_rom_0_freezer_io_in_rd),
    .io_in_addr(sound_io_rom_0_freezer_io_in_addr),
    .io_in_dout(sound_io_rom_0_freezer_io_in_dout),
    .io_in_wait_n(sound_io_rom_0_freezer_io_in_wait_n),
    .io_in_valid(sound_io_rom_0_freezer_io_in_valid),
    .io_out_rd(sound_io_rom_0_freezer_io_out_rd),
    .io_out_addr(sound_io_rom_0_freezer_io_out_addr),
    .io_out_dout(sound_io_rom_0_freezer_io_out_dout),
    .io_out_wait_n(sound_io_rom_0_freezer_io_out_wait_n),
    .io_out_valid(sound_io_rom_0_freezer_io_out_valid)
  );
  ReadDataFreezer_1 sound_io_rom_1_freezer ( // @[Crossing.scala 213:25]
    .clock(sound_io_rom_1_freezer_clock),
    .reset(sound_io_rom_1_freezer_reset),
    .io_targetClock(sound_io_rom_1_freezer_io_targetClock),
    .io_in_rd(sound_io_rom_1_freezer_io_in_rd),
    .io_in_addr(sound_io_rom_1_freezer_io_in_addr),
    .io_in_dout(sound_io_rom_1_freezer_io_in_dout),
    .io_in_wait_n(sound_io_rom_1_freezer_io_in_wait_n),
    .io_in_valid(sound_io_rom_1_freezer_io_in_valid),
    .io_out_rd(sound_io_rom_1_freezer_io_out_rd),
    .io_out_addr(sound_io_rom_1_freezer_io_out_addr),
    .io_out_dout(sound_io_rom_1_freezer_io_out_dout),
    .io_out_wait_n(sound_io_rom_1_freezer_io_out_wait_n),
    .io_out_valid(sound_io_rom_1_freezer_io_out_valid)
  );
  GPU gpu ( // @[Cave.scala 163:19]
    .clock(gpu_clock),
    .reset(gpu_reset),
    .io_videoClock(gpu_io_videoClock),
    .io_layerCtrl_0_enable(gpu_io_layerCtrl_0_enable),
    .io_layerCtrl_0_format(gpu_io_layerCtrl_0_format),
    .io_layerCtrl_0_regs_tileSize(gpu_io_layerCtrl_0_regs_tileSize),
    .io_layerCtrl_0_regs_enable(gpu_io_layerCtrl_0_regs_enable),
    .io_layerCtrl_0_regs_flipX(gpu_io_layerCtrl_0_regs_flipX),
    .io_layerCtrl_0_regs_flipY(gpu_io_layerCtrl_0_regs_flipY),
    .io_layerCtrl_0_regs_rowScrollEnable(gpu_io_layerCtrl_0_regs_rowScrollEnable),
    .io_layerCtrl_0_regs_rowSelectEnable(gpu_io_layerCtrl_0_regs_rowSelectEnable),
    .io_layerCtrl_0_regs_scroll_x(gpu_io_layerCtrl_0_regs_scroll_x),
    .io_layerCtrl_0_regs_scroll_y(gpu_io_layerCtrl_0_regs_scroll_y),
    .io_layerCtrl_0_vram8x8_addr(gpu_io_layerCtrl_0_vram8x8_addr),
    .io_layerCtrl_0_vram8x8_dout(gpu_io_layerCtrl_0_vram8x8_dout),
    .io_layerCtrl_0_vram16x16_addr(gpu_io_layerCtrl_0_vram16x16_addr),
    .io_layerCtrl_0_vram16x16_dout(gpu_io_layerCtrl_0_vram16x16_dout),
    .io_layerCtrl_0_lineRam_addr(gpu_io_layerCtrl_0_lineRam_addr),
    .io_layerCtrl_0_lineRam_dout(gpu_io_layerCtrl_0_lineRam_dout),
    .io_layerCtrl_0_tileRom_rd(gpu_io_layerCtrl_0_tileRom_rd),
    .io_layerCtrl_0_tileRom_addr(gpu_io_layerCtrl_0_tileRom_addr),
    .io_layerCtrl_0_tileRom_dout(gpu_io_layerCtrl_0_tileRom_dout),
    .io_layerCtrl_1_enable(gpu_io_layerCtrl_1_enable),
    .io_layerCtrl_1_format(gpu_io_layerCtrl_1_format),
    .io_layerCtrl_1_regs_tileSize(gpu_io_layerCtrl_1_regs_tileSize),
    .io_layerCtrl_1_regs_enable(gpu_io_layerCtrl_1_regs_enable),
    .io_layerCtrl_1_regs_flipX(gpu_io_layerCtrl_1_regs_flipX),
    .io_layerCtrl_1_regs_flipY(gpu_io_layerCtrl_1_regs_flipY),
    .io_layerCtrl_1_regs_rowScrollEnable(gpu_io_layerCtrl_1_regs_rowScrollEnable),
    .io_layerCtrl_1_regs_rowSelectEnable(gpu_io_layerCtrl_1_regs_rowSelectEnable),
    .io_layerCtrl_1_regs_scroll_x(gpu_io_layerCtrl_1_regs_scroll_x),
    .io_layerCtrl_1_regs_scroll_y(gpu_io_layerCtrl_1_regs_scroll_y),
    .io_layerCtrl_1_vram8x8_addr(gpu_io_layerCtrl_1_vram8x8_addr),
    .io_layerCtrl_1_vram8x8_dout(gpu_io_layerCtrl_1_vram8x8_dout),
    .io_layerCtrl_1_vram16x16_addr(gpu_io_layerCtrl_1_vram16x16_addr),
    .io_layerCtrl_1_vram16x16_dout(gpu_io_layerCtrl_1_vram16x16_dout),
    .io_layerCtrl_1_lineRam_addr(gpu_io_layerCtrl_1_lineRam_addr),
    .io_layerCtrl_1_lineRam_dout(gpu_io_layerCtrl_1_lineRam_dout),
    .io_layerCtrl_1_tileRom_rd(gpu_io_layerCtrl_1_tileRom_rd),
    .io_layerCtrl_1_tileRom_addr(gpu_io_layerCtrl_1_tileRom_addr),
    .io_layerCtrl_1_tileRom_dout(gpu_io_layerCtrl_1_tileRom_dout),
    .io_layerCtrl_2_enable(gpu_io_layerCtrl_2_enable),
    .io_layerCtrl_2_format(gpu_io_layerCtrl_2_format),
    .io_layerCtrl_2_regs_tileSize(gpu_io_layerCtrl_2_regs_tileSize),
    .io_layerCtrl_2_regs_enable(gpu_io_layerCtrl_2_regs_enable),
    .io_layerCtrl_2_regs_flipX(gpu_io_layerCtrl_2_regs_flipX),
    .io_layerCtrl_2_regs_flipY(gpu_io_layerCtrl_2_regs_flipY),
    .io_layerCtrl_2_regs_rowScrollEnable(gpu_io_layerCtrl_2_regs_rowScrollEnable),
    .io_layerCtrl_2_regs_rowSelectEnable(gpu_io_layerCtrl_2_regs_rowSelectEnable),
    .io_layerCtrl_2_regs_scroll_x(gpu_io_layerCtrl_2_regs_scroll_x),
    .io_layerCtrl_2_regs_scroll_y(gpu_io_layerCtrl_2_regs_scroll_y),
    .io_layerCtrl_2_vram8x8_addr(gpu_io_layerCtrl_2_vram8x8_addr),
    .io_layerCtrl_2_vram8x8_dout(gpu_io_layerCtrl_2_vram8x8_dout),
    .io_layerCtrl_2_vram16x16_addr(gpu_io_layerCtrl_2_vram16x16_addr),
    .io_layerCtrl_2_vram16x16_dout(gpu_io_layerCtrl_2_vram16x16_dout),
    .io_layerCtrl_2_lineRam_addr(gpu_io_layerCtrl_2_lineRam_addr),
    .io_layerCtrl_2_lineRam_dout(gpu_io_layerCtrl_2_lineRam_dout),
    .io_layerCtrl_2_tileRom_rd(gpu_io_layerCtrl_2_tileRom_rd),
    .io_layerCtrl_2_tileRom_addr(gpu_io_layerCtrl_2_tileRom_addr),
    .io_layerCtrl_2_tileRom_dout(gpu_io_layerCtrl_2_tileRom_dout),
    .io_spriteCtrl_enable(gpu_io_spriteCtrl_enable),
    .io_spriteCtrl_format(gpu_io_spriteCtrl_format),
    .io_spriteCtrl_start(gpu_io_spriteCtrl_start),
    .io_spriteCtrl_zoom(gpu_io_spriteCtrl_zoom),
    .io_spriteCtrl_regs_offset_x(gpu_io_spriteCtrl_regs_offset_x),
    .io_spriteCtrl_regs_offset_y(gpu_io_spriteCtrl_regs_offset_y),
    .io_spriteCtrl_regs_bank(gpu_io_spriteCtrl_regs_bank),
    .io_spriteCtrl_regs_fixed(gpu_io_spriteCtrl_regs_fixed),
    .io_spriteCtrl_regs_hFlip(gpu_io_spriteCtrl_regs_hFlip),
    .io_spriteCtrl_vram_rd(gpu_io_spriteCtrl_vram_rd),
    .io_spriteCtrl_vram_addr(gpu_io_spriteCtrl_vram_addr),
    .io_spriteCtrl_vram_dout(gpu_io_spriteCtrl_vram_dout),
    .io_spriteCtrl_tileRom_rd(gpu_io_spriteCtrl_tileRom_rd),
    .io_spriteCtrl_tileRom_addr(gpu_io_spriteCtrl_tileRom_addr),
    .io_spriteCtrl_tileRom_dout(gpu_io_spriteCtrl_tileRom_dout),
    .io_spriteCtrl_tileRom_wait_n(gpu_io_spriteCtrl_tileRom_wait_n),
    .io_spriteCtrl_tileRom_valid(gpu_io_spriteCtrl_tileRom_valid),
    .io_spriteCtrl_tileRom_burstLength(gpu_io_spriteCtrl_tileRom_burstLength),
    .io_spriteCtrl_tileRom_burstDone(gpu_io_spriteCtrl_tileRom_burstDone),
    .io_gameConfig_granularity(gpu_io_gameConfig_granularity),
    .io_gameConfig_layer_0_paletteBank(gpu_io_gameConfig_layer_0_paletteBank),
    .io_gameConfig_layer_1_paletteBank(gpu_io_gameConfig_layer_1_paletteBank),
    .io_gameConfig_layer_2_paletteBank(gpu_io_gameConfig_layer_2_paletteBank),
    .io_options_rotate(gpu_io_options_rotate),
    .io_options_flip(gpu_io_options_flip),
    .io_video_clockEnable(gpu_io_video_clockEnable),
    .io_video_displayEnable(gpu_io_video_displayEnable),
    .io_video_pos_x(gpu_io_video_pos_x),
    .io_video_pos_y(gpu_io_video_pos_y),
    .io_video_vBlank(gpu_io_video_vBlank),
    .io_video_regs_size_x(gpu_io_video_regs_size_x),
    .io_video_regs_size_y(gpu_io_video_regs_size_y),
    .io_spriteLineBuffer_addr(gpu_io_spriteLineBuffer_addr),
    .io_spriteLineBuffer_dout(gpu_io_spriteLineBuffer_dout),
    .io_spriteFrameBuffer_wr(gpu_io_spriteFrameBuffer_wr),
    .io_spriteFrameBuffer_addr(gpu_io_spriteFrameBuffer_addr),
    .io_spriteFrameBuffer_din(gpu_io_spriteFrameBuffer_din),
    .io_spriteFrameBuffer_wait_n(gpu_io_spriteFrameBuffer_wait_n),
    .io_systemFrameBuffer_wr(gpu_io_systemFrameBuffer_wr),
    .io_systemFrameBuffer_addr(gpu_io_systemFrameBuffer_addr),
    .io_systemFrameBuffer_din(gpu_io_systemFrameBuffer_din),
    .io_paletteRam_addr(gpu_io_paletteRam_addr),
    .io_paletteRam_dout(gpu_io_paletteRam_dout),
    .io_rgb(gpu_io_rgb)
  );
  Crossing gpu_io_layerCtrl_0_tileRom_crossing ( // @[Crossing.scala 200:26]
    .clock(gpu_io_layerCtrl_0_tileRom_crossing_clock),
    .io_targetClock(gpu_io_layerCtrl_0_tileRom_crossing_io_targetClock),
    .io_in_rd(gpu_io_layerCtrl_0_tileRom_crossing_io_in_rd),
    .io_in_addr(gpu_io_layerCtrl_0_tileRom_crossing_io_in_addr),
    .io_in_dout(gpu_io_layerCtrl_0_tileRom_crossing_io_in_dout),
    .io_out_rd(gpu_io_layerCtrl_0_tileRom_crossing_io_out_rd),
    .io_out_addr(gpu_io_layerCtrl_0_tileRom_crossing_io_out_addr),
    .io_out_dout(gpu_io_layerCtrl_0_tileRom_crossing_io_out_dout),
    .io_out_wait_n(gpu_io_layerCtrl_0_tileRom_crossing_io_out_wait_n),
    .io_out_valid(gpu_io_layerCtrl_0_tileRom_crossing_io_out_valid)
  );
  Crossing gpu_io_layerCtrl_1_tileRom_crossing ( // @[Crossing.scala 200:26]
    .clock(gpu_io_layerCtrl_1_tileRom_crossing_clock),
    .io_targetClock(gpu_io_layerCtrl_1_tileRom_crossing_io_targetClock),
    .io_in_rd(gpu_io_layerCtrl_1_tileRom_crossing_io_in_rd),
    .io_in_addr(gpu_io_layerCtrl_1_tileRom_crossing_io_in_addr),
    .io_in_dout(gpu_io_layerCtrl_1_tileRom_crossing_io_in_dout),
    .io_out_rd(gpu_io_layerCtrl_1_tileRom_crossing_io_out_rd),
    .io_out_addr(gpu_io_layerCtrl_1_tileRom_crossing_io_out_addr),
    .io_out_dout(gpu_io_layerCtrl_1_tileRom_crossing_io_out_dout),
    .io_out_wait_n(gpu_io_layerCtrl_1_tileRom_crossing_io_out_wait_n),
    .io_out_valid(gpu_io_layerCtrl_1_tileRom_crossing_io_out_valid)
  );
  Crossing gpu_io_layerCtrl_2_tileRom_crossing ( // @[Crossing.scala 200:26]
    .clock(gpu_io_layerCtrl_2_tileRom_crossing_clock),
    .io_targetClock(gpu_io_layerCtrl_2_tileRom_crossing_io_targetClock),
    .io_in_rd(gpu_io_layerCtrl_2_tileRom_crossing_io_in_rd),
    .io_in_addr(gpu_io_layerCtrl_2_tileRom_crossing_io_in_addr),
    .io_in_dout(gpu_io_layerCtrl_2_tileRom_crossing_io_in_dout),
    .io_out_rd(gpu_io_layerCtrl_2_tileRom_crossing_io_out_rd),
    .io_out_addr(gpu_io_layerCtrl_2_tileRom_crossing_io_out_addr),
    .io_out_dout(gpu_io_layerCtrl_2_tileRom_crossing_io_out_dout),
    .io_out_wait_n(gpu_io_layerCtrl_2_tileRom_crossing_io_out_wait_n),
    .io_out_valid(gpu_io_layerCtrl_2_tileRom_crossing_io_out_valid)
  );
  SpriteFrameBuffer spriteFrameBuffer ( // @[Cave.scala 187:33]
    .clock(spriteFrameBuffer_clock),
    .reset(spriteFrameBuffer_reset),
    .io_videoClock(spriteFrameBuffer_io_videoClock),
    .io_enable(spriteFrameBuffer_io_enable),
    .io_swap(spriteFrameBuffer_io_swap),
    .io_video_pos_y(spriteFrameBuffer_io_video_pos_y),
    .io_video_hBlank(spriteFrameBuffer_io_video_hBlank),
    .io_lineBuffer_addr(spriteFrameBuffer_io_lineBuffer_addr),
    .io_lineBuffer_dout(spriteFrameBuffer_io_lineBuffer_dout),
    .io_frameBuffer_wr(spriteFrameBuffer_io_frameBuffer_wr),
    .io_frameBuffer_addr(spriteFrameBuffer_io_frameBuffer_addr),
    .io_frameBuffer_din(spriteFrameBuffer_io_frameBuffer_din),
    .io_frameBuffer_wait_n(spriteFrameBuffer_io_frameBuffer_wait_n),
    .io_ddr_rd(spriteFrameBuffer_io_ddr_rd),
    .io_ddr_wr(spriteFrameBuffer_io_ddr_wr),
    .io_ddr_addr(spriteFrameBuffer_io_ddr_addr),
    .io_ddr_mask(spriteFrameBuffer_io_ddr_mask),
    .io_ddr_din(spriteFrameBuffer_io_ddr_din),
    .io_ddr_dout(spriteFrameBuffer_io_ddr_dout),
    .io_ddr_wait_n(spriteFrameBuffer_io_ddr_wait_n),
    .io_ddr_valid(spriteFrameBuffer_io_ddr_valid),
    .io_ddr_burstLength(spriteFrameBuffer_io_ddr_burstLength),
    .io_ddr_burstDone(spriteFrameBuffer_io_ddr_burstDone)
  );
  SystemFrameBuffer systemFrameBuffer ( // @[Cave.scala 197:33]
    .clock(systemFrameBuffer_clock),
    .reset(systemFrameBuffer_reset),
    .io_videoClock(systemFrameBuffer_io_videoClock),
    .io_enable(systemFrameBuffer_io_enable),
    .io_rotate(systemFrameBuffer_io_rotate),
    .io_forceBlank(systemFrameBuffer_io_forceBlank),
    .io_video_vBlank(systemFrameBuffer_io_video_vBlank),
    .io_video_regs_size_x(systemFrameBuffer_io_video_regs_size_x),
    .io_video_regs_size_y(systemFrameBuffer_io_video_regs_size_y),
    .io_frameBufferCtrl_enable(systemFrameBuffer_io_frameBufferCtrl_enable),
    .io_frameBufferCtrl_hSize(systemFrameBuffer_io_frameBufferCtrl_hSize),
    .io_frameBufferCtrl_vSize(systemFrameBuffer_io_frameBufferCtrl_vSize),
    .io_frameBufferCtrl_baseAddr(systemFrameBuffer_io_frameBufferCtrl_baseAddr),
    .io_frameBufferCtrl_stride(systemFrameBuffer_io_frameBufferCtrl_stride),
    .io_frameBufferCtrl_vBlank(systemFrameBuffer_io_frameBufferCtrl_vBlank),
    .io_frameBufferCtrl_lowLat(systemFrameBuffer_io_frameBufferCtrl_lowLat),
    .io_frameBufferCtrl_forceBlank(systemFrameBuffer_io_frameBufferCtrl_forceBlank),
    .io_frameBuffer_wr(systemFrameBuffer_io_frameBuffer_wr),
    .io_frameBuffer_addr(systemFrameBuffer_io_frameBuffer_addr),
    .io_frameBuffer_din(systemFrameBuffer_io_frameBuffer_din),
    .io_ddr_wr(systemFrameBuffer_io_ddr_wr),
    .io_ddr_addr(systemFrameBuffer_io_ddr_addr),
    .io_ddr_mask(systemFrameBuffer_io_ddr_mask),
    .io_ddr_din(systemFrameBuffer_io_ddr_din),
    .io_ddr_wait_n(systemFrameBuffer_io_ddr_wait_n)
  );
  assign ioctl_wait_n = videoSys_io_prog_video_writeEnable | _GEN_8; // @[IOCTL.scala 109:{23,32}]
  assign ioctl_din = memSys_io_prog_nvram_readEnable ? memSys_io_prog_nvram_view__ioctl_din_r : 16'h0; // @[IOCTL.scala 88:{22,28} 62:9]
  assign led_power = 1'h0; // @[Cave.scala 211:16]
  assign led_disk = ioctl_download; // @[Cave.scala 212:15]
  assign led_user = memSys_io_ready; // @[Cave.scala 213:15]
  assign frameBufferCtrl_enable = systemFrameBuffer_io_frameBufferCtrl_enable; // @[Cave.scala 203:40]
  assign frameBufferCtrl_hSize = systemFrameBuffer_io_frameBufferCtrl_hSize; // @[Cave.scala 203:40]
  assign frameBufferCtrl_vSize = systemFrameBuffer_io_frameBufferCtrl_vSize; // @[Cave.scala 203:40]
  assign frameBufferCtrl_format = 5'h6; // @[Cave.scala 203:40]
  assign frameBufferCtrl_baseAddr = systemFrameBuffer_io_frameBufferCtrl_baseAddr; // @[Cave.scala 203:40]
  assign frameBufferCtrl_stride = systemFrameBuffer_io_frameBufferCtrl_stride; // @[Cave.scala 203:40]
  assign frameBufferCtrl_forceBlank = systemFrameBuffer_io_frameBufferCtrl_forceBlank; // @[Cave.scala 203:40]
  assign video_clockEnable = videoSys_io_video_clockEnable; // @[Cave.scala 208:12]
  assign video_displayEnable = videoSys_io_video_displayEnable; // @[Cave.scala 208:12]
  assign video_pos_x = videoSys_io_video_pos_x; // @[Cave.scala 208:12]
  assign video_pos_y = videoSys_io_video_pos_y; // @[Cave.scala 208:12]
  assign video_hSync = videoSys_io_video_hSync; // @[Cave.scala 208:12]
  assign video_vSync = videoSys_io_video_vSync; // @[Cave.scala 208:12]
  assign video_hBlank = videoSys_io_video_hBlank; // @[Cave.scala 208:12]
  assign video_vBlank = videoSys_io_video_vBlank; // @[Cave.scala 208:12]
  assign video_regs_size_x = videoSys_io_video_regs_size_x; // @[Cave.scala 208:12]
  assign video_regs_size_y = videoSys_io_video_regs_size_y; // @[Cave.scala 208:12]
  assign video_regs_frontPorch_x = videoSys_io_video_regs_frontPorch_x; // @[Cave.scala 208:12]
  assign video_regs_frontPorch_y = videoSys_io_video_regs_frontPorch_y; // @[Cave.scala 208:12]
  assign video_regs_retrace_x = videoSys_io_video_regs_retrace_x; // @[Cave.scala 208:12]
  assign video_regs_retrace_y = videoSys_io_video_regs_retrace_y; // @[Cave.scala 208:12]
  assign video_changeMode = videoSys_io_video_changeMode; // @[Cave.scala 208:12]
  assign rgb = gpu_io_rgb; // @[Cave.scala 209:10]
  assign audio = sound_io_audio; // @[Cave.scala 210:12]
  assign sdram_cke = 1'h1; // @[Cave.scala 123:18]
  assign sdram_cs_n = sdram_1_io_sdram_cs_n; // @[Cave.scala 123:18]
  assign sdram_ras_n = sdram_1_io_sdram_ras_n; // @[Cave.scala 123:18]
  assign sdram_cas_n = sdram_1_io_sdram_cas_n; // @[Cave.scala 123:18]
  assign sdram_we_n = sdram_1_io_sdram_we_n; // @[Cave.scala 123:18]
  assign sdram_oe_n = sdram_1_io_sdram_oe_n; // @[Cave.scala 123:18]
  assign sdram_bank = sdram_1_io_sdram_bank; // @[Cave.scala 123:18]
  assign sdram_addr = sdram_1_io_sdram_addr; // @[Cave.scala 123:18]
  assign sdram_din = sdram_1_io_sdram_din; // @[Cave.scala 123:18]
  assign ddr_rd = ddr_1_io_ddr_rd; // @[Cave.scala 119:14]
  assign ddr_wr = ddr_1_io_ddr_wr; // @[Cave.scala 119:14]
  assign ddr_addr = ddr_1_io_ddr_addr; // @[Cave.scala 119:14]
  assign ddr_mask = ddr_1_io_ddr_mask; // @[Cave.scala 119:14]
  assign ddr_din = ddr_1_io_ddr_din; // @[Cave.scala 119:14]
  assign ddr_burstLength = ddr_1_io_ddr_burstLength; // @[Cave.scala 119:14]
  assign dipsRegs_clock = clock;
  assign dipsRegs_io_mem_wr = dipsRegs_io_mem_writeEnable & ioctl_wr; // @[IOCTL.scala 96:27]
  assign dipsRegs_io_mem_addr = ioctl_addr[2:1]; // @[Cave.scala 113:19]
  assign dipsRegs_io_mem_din = ioctl_dout; // @[IOCTL.scala 100:13 95:19]
  assign ddr_1_clock = clock;
  assign ddr_1_reset = reset;
  assign ddr_1_io_mem_rd = memSys_io_ddr_rd; // @[Cave.scala 131:17]
  assign ddr_1_io_mem_wr = memSys_io_ddr_wr; // @[Cave.scala 131:17]
  assign ddr_1_io_mem_addr = memSys_io_ddr_addr; // @[Cave.scala 131:17]
  assign ddr_1_io_mem_mask = memSys_io_ddr_mask; // @[Cave.scala 131:17]
  assign ddr_1_io_mem_din = memSys_io_ddr_din; // @[Cave.scala 131:17]
  assign ddr_1_io_mem_burstLength = memSys_io_ddr_burstLength; // @[Cave.scala 131:17]
  assign ddr_1_io_ddr_dout = ddr_dout; // @[Cave.scala 119:14]
  assign ddr_1_io_ddr_wait_n = ddr_wait_n; // @[Cave.scala 119:14]
  assign ddr_1_io_ddr_valid = ddr_valid; // @[Cave.scala 119:14]
  assign sdram_1_clock = clock;
  assign sdram_1_reset = reset;
  assign sdram_1_io_mem_rd = memSys_io_sdram_rd; // @[Cave.scala 132:19]
  assign sdram_1_io_mem_wr = memSys_io_sdram_wr; // @[Cave.scala 132:19]
  assign sdram_1_io_mem_addr = memSys_io_sdram_addr; // @[Cave.scala 132:19]
  assign sdram_1_io_mem_din = memSys_io_sdram_din; // @[Cave.scala 132:19]
  assign sdram_1_io_sdram_dout = sdram_dout; // @[Cave.scala 123:18]
  assign memSys_clock = clock;
  assign memSys_reset = reset;
  assign memSys_io_gameConfig_eepromOffset = 4'h4 == gameIndexReg ? 32'h100000 : _gameConfig_T_11_eepromOffset; // @[Mux.scala 81:58]
  assign memSys_io_gameConfig_sound_0_romOffset = 4'h4 == gameIndexReg ? 32'h100080 : _gameConfig_T_11_sound_0_romOffset
    ; // @[Mux.scala 81:58]
  assign memSys_io_gameConfig_sound_1_romOffset = 4'h4 == gameIndexReg ? 32'h0 : _gameConfig_T_11_sound_1_romOffset; // @[Mux.scala 81:58]
  assign memSys_io_gameConfig_layer_0_romOffset = 4'h4 == gameIndexReg ? 32'h300080 : _gameConfig_T_11_layer_0_romOffset
    ; // @[Mux.scala 81:58]
  assign memSys_io_gameConfig_layer_1_romOffset = 4'h4 == gameIndexReg ? 32'h0 : _gameConfig_T_11_layer_1_romOffset; // @[Mux.scala 81:58]
  assign memSys_io_gameConfig_layer_2_romOffset = 4'h4 == gameIndexReg ? 32'h0 : _gameConfig_T_11_layer_2_romOffset; // @[Mux.scala 81:58]
  assign memSys_io_gameConfig_sprite_romOffset = 4'h4 == gameIndexReg ? 32'h700080 : _gameConfig_T_11_sprite_romOffset; // @[Mux.scala 81:58]
  assign memSys_io_prog_rom_wr = memSys_io_prog_rom_writeEnable & ioctl_wr; // @[IOCTL.scala 69:27]
  assign memSys_io_prog_rom_addr = ioctl_addr; // @[IOCTL.scala 68:19 71:14]
  assign memSys_io_prog_rom_din = ioctl_dout; // @[IOCTL.scala 68:19 73:13]
  assign memSys_io_prog_nvram_rd = memSys_io_prog_nvram_readEnable & ioctl_rd; // @[IOCTL.scala 82:26]
  assign memSys_io_prog_nvram_wr = memSys_io_prog_nvram_writeEnable & ioctl_wr; // @[IOCTL.scala 83:27]
  assign memSys_io_prog_nvram_addr = ioctl_addr; // @[IOCTL.scala 81:19 85:14]
  assign memSys_io_prog_nvram_din = ioctl_dout; // @[IOCTL.scala 81:19 87:13]
  assign memSys_io_prog_done = _memSys_io_prog_done_T_1 & _memSys_io_prog_rom_writeEnable_T; // @[Cave.scala 130:58]
  assign memSys_io_progRom_rd = main_io_progRom_freezer_io_out_rd; // @[Crossing.scala 215:20]
  assign memSys_io_progRom_addr = main_io_progRom_freezer_io_out_addr; // @[Crossing.scala 215:20]
  assign memSys_io_eeprom_rd = main_io_eeprom_freezer_io_out_rd; // @[Crossing.scala 228:20]
  assign memSys_io_eeprom_wr = main_io_eeprom_freezer_io_out_wr; // @[Crossing.scala 228:20]
  assign memSys_io_eeprom_addr = main_io_eeprom_freezer_io_out_addr; // @[Crossing.scala 228:20]
  assign memSys_io_eeprom_din = main_io_eeprom_freezer_io_out_din; // @[Crossing.scala 228:20]
  assign memSys_io_soundRom_0_rd = sound_io_rom_0_freezer_io_out_rd; // @[Crossing.scala 215:20]
  assign memSys_io_soundRom_0_addr = sound_io_rom_0_freezer_io_out_addr; // @[Crossing.scala 215:20]
  assign memSys_io_soundRom_1_rd = sound_io_rom_1_freezer_io_out_rd; // @[Crossing.scala 215:20]
  assign memSys_io_soundRom_1_addr = sound_io_rom_1_freezer_io_out_addr; // @[Crossing.scala 215:20]
  assign memSys_io_layerTileRom_0_rd = gpu_io_layerCtrl_0_tileRom_crossing_io_out_rd; // @[Crossing.scala 202:21]
  assign memSys_io_layerTileRom_0_addr = gpu_io_layerCtrl_0_tileRom_crossing_io_out_addr; // @[Crossing.scala 202:21]
  assign memSys_io_layerTileRom_1_rd = gpu_io_layerCtrl_1_tileRom_crossing_io_out_rd; // @[Crossing.scala 202:21]
  assign memSys_io_layerTileRom_1_addr = gpu_io_layerCtrl_1_tileRom_crossing_io_out_addr; // @[Crossing.scala 202:21]
  assign memSys_io_layerTileRom_2_rd = gpu_io_layerCtrl_2_tileRom_crossing_io_out_rd; // @[Crossing.scala 202:21]
  assign memSys_io_layerTileRom_2_addr = gpu_io_layerCtrl_2_tileRom_crossing_io_out_addr; // @[Crossing.scala 202:21]
  assign memSys_io_spriteTileRom_rd = gpu_io_spriteCtrl_tileRom_rd; // @[Cave.scala 179:29]
  assign memSys_io_spriteTileRom_addr = gpu_io_spriteCtrl_tileRom_addr; // @[Cave.scala 179:29]
  assign memSys_io_spriteTileRom_burstLength = gpu_io_spriteCtrl_tileRom_burstLength; // @[Cave.scala 179:29]
  assign memSys_io_ddr_dout = ddr_1_io_mem_dout; // @[Cave.scala 131:17]
  assign memSys_io_ddr_wait_n = ddr_1_io_mem_wait_n; // @[Cave.scala 131:17]
  assign memSys_io_ddr_valid = ddr_1_io_mem_valid; // @[Cave.scala 131:17]
  assign memSys_io_ddr_burstDone = ddr_1_io_mem_burstDone; // @[Cave.scala 131:17]
  assign memSys_io_sdram_dout = sdram_1_io_mem_dout; // @[Cave.scala 132:19]
  assign memSys_io_sdram_wait_n = sdram_1_io_mem_wait_n; // @[Cave.scala 132:19]
  assign memSys_io_sdram_valid = sdram_1_io_mem_valid; // @[Cave.scala 132:19]
  assign memSys_io_sdram_burstDone = sdram_1_io_mem_burstDone; // @[Cave.scala 132:19]
  assign memSys_io_spriteFrameBuffer_rd = spriteFrameBuffer_io_ddr_rd; // @[Cave.scala 194:28]
  assign memSys_io_spriteFrameBuffer_wr = spriteFrameBuffer_io_ddr_wr; // @[Cave.scala 194:28]
  assign memSys_io_spriteFrameBuffer_addr = spriteFrameBuffer_io_ddr_addr; // @[Cave.scala 194:28]
  assign memSys_io_spriteFrameBuffer_mask = spriteFrameBuffer_io_ddr_mask; // @[Cave.scala 194:28]
  assign memSys_io_spriteFrameBuffer_din = spriteFrameBuffer_io_ddr_din; // @[Cave.scala 194:28]
  assign memSys_io_spriteFrameBuffer_burstLength = spriteFrameBuffer_io_ddr_burstLength; // @[Cave.scala 194:28]
  assign memSys_io_systemFrameBuffer_wr = systemFrameBuffer_io_ddr_wr; // @[Cave.scala 205:28]
  assign memSys_io_systemFrameBuffer_addr = systemFrameBuffer_io_ddr_addr; // @[Cave.scala 205:28]
  assign memSys_io_systemFrameBuffer_mask = systemFrameBuffer_io_ddr_mask; // @[Cave.scala 205:28]
  assign memSys_io_systemFrameBuffer_din = systemFrameBuffer_io_ddr_din; // @[Cave.scala 205:28]
  assign videoSys_clock = clock;
  assign videoSys_reset = reset;
  assign videoSys_io_videoClock = videoClock; // @[Cave.scala 136:26]
  assign videoSys_io_videoReset = videoReset; // @[Cave.scala 137:26]
  assign videoSys_io_prog_video_wr = videoSys_io_prog_video_writeEnable & ioctl_wr; // @[IOCTL.scala 108:27]
  assign videoSys_io_prog_video_addr = ioctl_addr; // @[IOCTL.scala 107:19 110:14]
  assign videoSys_io_prog_video_din = ioctl_dout; // @[IOCTL.scala 107:19 112:13]
  assign videoSys_io_prog_done = _videoSys_io_prog_done_T_1 & _videoSys_io_prog_video_writeEnable_T; // @[Cave.scala 139:60]
  assign videoSys_io_options_offset_x = options_offset_x; // @[Cave.scala 140:23]
  assign videoSys_io_options_offset_y = options_offset_y; // @[Cave.scala 140:23]
  assign videoSys_io_options_compatibility = options_compatibility; // @[Cave.scala 140:23]
  assign main_clock = cpuClock;
  assign main_reset = cpuReset | ~memSys_io_ready; // @[Cave.scala 143:57]
  assign main_io_videoClock = videoClock; // @[Cave.scala 144:22]
  assign main_io_spriteClock = clock; // @[Cave.scala 145:23]
  assign main_io_gameIndex = gameIndexReg; // @[Cave.scala 146:21]
  assign main_io_options_service = options_service; // @[Cave.scala 147:19]
  assign main_io_player_0_up = player_0_up; // @[Cave.scala 149:18]
  assign main_io_player_0_down = player_0_down; // @[Cave.scala 149:18]
  assign main_io_player_0_left = player_0_left; // @[Cave.scala 149:18]
  assign main_io_player_0_right = player_0_right; // @[Cave.scala 149:18]
  assign main_io_player_0_buttons = player_0_buttons; // @[Cave.scala 149:18]
  assign main_io_player_0_start = player_0_start; // @[Cave.scala 149:18]
  assign main_io_player_0_coin = player_0_coin; // @[Cave.scala 149:18]
  assign main_io_player_0_pause = player_0_pause; // @[Cave.scala 149:18]
  assign main_io_player_1_up = player_1_up; // @[Cave.scala 149:18]
  assign main_io_player_1_down = player_1_down; // @[Cave.scala 149:18]
  assign main_io_player_1_left = player_1_left; // @[Cave.scala 149:18]
  assign main_io_player_1_right = player_1_right; // @[Cave.scala 149:18]
  assign main_io_player_1_buttons = player_1_buttons; // @[Cave.scala 149:18]
  assign main_io_player_1_start = player_1_start; // @[Cave.scala 149:18]
  assign main_io_player_1_coin = player_1_coin; // @[Cave.scala 149:18]
  assign main_io_player_1_pause = player_1_pause; // @[Cave.scala 149:18]
  assign main_io_dips_0 = dipsRegs_io_regs_0; // @[Cave.scala 148:16]
  assign main_io_video_vBlank = videoSys_io_video_vBlank; // @[Cave.scala 150:17]
  assign main_io_gpuMem_layer_0_vram8x8_addr = gpu_io_layerCtrl_0_vram8x8_addr; // @[Cave.scala 168:33]
  assign main_io_gpuMem_layer_0_vram16x16_addr = gpu_io_layerCtrl_0_vram16x16_addr; // @[Cave.scala 169:35]
  assign main_io_gpuMem_layer_0_lineRam_addr = gpu_io_layerCtrl_0_lineRam_addr; // @[Cave.scala 170:33]
  assign main_io_gpuMem_layer_1_vram8x8_addr = gpu_io_layerCtrl_1_vram8x8_addr; // @[Cave.scala 168:33]
  assign main_io_gpuMem_layer_1_vram16x16_addr = gpu_io_layerCtrl_1_vram16x16_addr; // @[Cave.scala 169:35]
  assign main_io_gpuMem_layer_1_lineRam_addr = gpu_io_layerCtrl_1_lineRam_addr; // @[Cave.scala 170:33]
  assign main_io_gpuMem_layer_2_vram8x8_addr = gpu_io_layerCtrl_2_vram8x8_addr; // @[Cave.scala 168:33]
  assign main_io_gpuMem_layer_2_vram16x16_addr = gpu_io_layerCtrl_2_vram16x16_addr; // @[Cave.scala 169:35]
  assign main_io_gpuMem_layer_2_lineRam_addr = gpu_io_layerCtrl_2_lineRam_addr; // @[Cave.scala 170:33]
  assign main_io_gpuMem_sprite_vram_rd = gpu_io_spriteCtrl_vram_rd; // @[Cave.scala 178:26]
  assign main_io_gpuMem_sprite_vram_addr = gpu_io_spriteCtrl_vram_addr; // @[Cave.scala 178:26]
  assign main_io_gpuMem_paletteRam_addr = gpu_io_paletteRam_addr; // @[Cave.scala 184:21]
  assign main_io_soundCtrl_oki_0_dout = sound_io_ctrl_oki_0_dout; // @[Cave.scala 158:17]
  assign main_io_soundCtrl_oki_1_dout = sound_io_ctrl_oki_1_dout; // @[Cave.scala 158:17]
  assign main_io_soundCtrl_ymz_dout = sound_io_ctrl_ymz_dout; // @[Cave.scala 158:17]
  assign main_io_soundCtrl_irq = sound_io_ctrl_irq; // @[Cave.scala 158:17]
  assign main_io_progRom_dout = main_io_progRom_freezer_io_in_dout; // @[Cave.scala 151:19]
  assign main_io_progRom_valid = main_io_progRom_freezer_io_in_valid; // @[Cave.scala 151:19]
  assign main_io_eeprom_dout = main_io_eeprom_freezer_io_in_dout; // @[Cave.scala 152:18]
  assign main_io_eeprom_wait_n = main_io_eeprom_freezer_io_in_wait_n; // @[Cave.scala 152:18]
  assign main_io_eeprom_valid = main_io_eeprom_freezer_io_in_valid; // @[Cave.scala 152:18]
  assign main_io_progRom_freezer_clock = clock;
  assign main_io_progRom_freezer_reset = reset;
  assign main_io_progRom_freezer_io_targetClock = cpuClock; // @[Crossing.scala 214:28]
  assign main_io_progRom_freezer_io_in_rd = main_io_progRom_rd; // @[Cave.scala 151:19]
  assign main_io_progRom_freezer_io_in_addr = main_io_progRom_addr; // @[Cave.scala 151:19]
  assign main_io_progRom_freezer_io_out_dout = memSys_io_progRom_dout; // @[Crossing.scala 215:20]
  assign main_io_progRom_freezer_io_out_wait_n = memSys_io_progRom_wait_n; // @[Crossing.scala 215:20]
  assign main_io_progRom_freezer_io_out_valid = memSys_io_progRom_valid; // @[Crossing.scala 215:20]
  assign main_io_eeprom_freezer_clock = clock;
  assign main_io_eeprom_freezer_reset = reset;
  assign main_io_eeprom_freezer_io_targetClock = cpuClock; // @[Crossing.scala 227:28]
  assign main_io_eeprom_freezer_io_in_rd = main_io_eeprom_rd; // @[Cave.scala 152:18]
  assign main_io_eeprom_freezer_io_in_wr = main_io_eeprom_wr; // @[Cave.scala 152:18]
  assign main_io_eeprom_freezer_io_in_addr = main_io_eeprom_addr; // @[Cave.scala 152:18]
  assign main_io_eeprom_freezer_io_in_din = main_io_eeprom_din; // @[Cave.scala 152:18]
  assign main_io_eeprom_freezer_io_out_dout = memSys_io_eeprom_dout; // @[Crossing.scala 228:20]
  assign main_io_eeprom_freezer_io_out_wait_n = memSys_io_eeprom_wait_n; // @[Crossing.scala 228:20]
  assign main_io_eeprom_freezer_io_out_valid = memSys_io_eeprom_valid; // @[Crossing.scala 228:20]
  assign sound_clock = cpuClock;
  assign sound_reset = cpuReset | _T; // @[Cave.scala 155:58]
  assign sound_io_ctrl_oki_0_wr = main_io_soundCtrl_oki_0_wr; // @[Cave.scala 158:17]
  assign sound_io_ctrl_oki_0_din = main_io_soundCtrl_oki_0_din; // @[Cave.scala 158:17]
  assign sound_io_ctrl_oki_1_wr = main_io_soundCtrl_oki_1_wr; // @[Cave.scala 158:17]
  assign sound_io_ctrl_oki_1_din = main_io_soundCtrl_oki_1_din; // @[Cave.scala 158:17]
  assign sound_io_ctrl_nmk_wr = main_io_soundCtrl_nmk_wr; // @[Cave.scala 158:17]
  assign sound_io_ctrl_nmk_addr = main_io_soundCtrl_nmk_addr; // @[Cave.scala 158:17]
  assign sound_io_ctrl_nmk_din = main_io_soundCtrl_nmk_din; // @[Cave.scala 158:17]
  assign sound_io_ctrl_ymz_rd = main_io_soundCtrl_ymz_rd; // @[Cave.scala 158:17]
  assign sound_io_ctrl_ymz_wr = main_io_soundCtrl_ymz_wr; // @[Cave.scala 158:17]
  assign sound_io_ctrl_ymz_addr = main_io_soundCtrl_ymz_addr; // @[Cave.scala 158:17]
  assign sound_io_ctrl_ymz_din = main_io_soundCtrl_ymz_din; // @[Cave.scala 158:17]
  assign sound_io_ctrl_req = main_io_soundCtrl_req; // @[Cave.scala 158:17]
  assign sound_io_ctrl_data = main_io_soundCtrl_data; // @[Cave.scala 158:17]
  assign sound_io_gameIndex = gameIndexReg; // @[Cave.scala 156:22]
  assign sound_io_gameConfig_sound_0_device = 4'h4 == gameIndexReg ? 2'h1 : _gameConfig_T_11_sound_0_device; // @[Mux.scala 81:58]
  assign sound_io_rom_0_dout = sound_io_rom_0_freezer_io_in_dout; // @[Cave.scala 159:19]
  assign sound_io_rom_0_wait_n = sound_io_rom_0_freezer_io_in_wait_n; // @[Cave.scala 159:19]
  assign sound_io_rom_0_valid = sound_io_rom_0_freezer_io_in_valid; // @[Cave.scala 159:19]
  assign sound_io_rom_1_dout = sound_io_rom_1_freezer_io_in_dout; // @[Cave.scala 160:19]
  assign sound_io_rom_1_valid = sound_io_rom_1_freezer_io_in_valid; // @[Cave.scala 160:19]
  assign sound_io_rom_0_freezer_clock = clock;
  assign sound_io_rom_0_freezer_reset = reset;
  assign sound_io_rom_0_freezer_io_targetClock = cpuClock; // @[Crossing.scala 214:28]
  assign sound_io_rom_0_freezer_io_in_rd = sound_io_rom_0_rd; // @[Cave.scala 159:19]
  assign sound_io_rom_0_freezer_io_in_addr = sound_io_rom_0_addr; // @[Cave.scala 159:19]
  assign sound_io_rom_0_freezer_io_out_dout = memSys_io_soundRom_0_dout; // @[Crossing.scala 215:20]
  assign sound_io_rom_0_freezer_io_out_wait_n = memSys_io_soundRom_0_wait_n; // @[Crossing.scala 215:20]
  assign sound_io_rom_0_freezer_io_out_valid = memSys_io_soundRom_0_valid; // @[Crossing.scala 215:20]
  assign sound_io_rom_1_freezer_clock = clock;
  assign sound_io_rom_1_freezer_reset = reset;
  assign sound_io_rom_1_freezer_io_targetClock = cpuClock; // @[Crossing.scala 214:28]
  assign sound_io_rom_1_freezer_io_in_rd = 1'h1; // @[Cave.scala 160:19]
  assign sound_io_rom_1_freezer_io_in_addr = sound_io_rom_1_addr; // @[Cave.scala 160:19]
  assign sound_io_rom_1_freezer_io_out_dout = memSys_io_soundRom_1_dout; // @[Crossing.scala 215:20]
  assign sound_io_rom_1_freezer_io_out_wait_n = memSys_io_soundRom_1_wait_n; // @[Crossing.scala 215:20]
  assign sound_io_rom_1_freezer_io_out_valid = memSys_io_soundRom_1_valid; // @[Crossing.scala 215:20]
  assign gpu_clock = clock;
  assign gpu_reset = reset;
  assign gpu_io_videoClock = videoClock; // @[Cave.scala 164:21]
  assign gpu_io_layerCtrl_0_enable = options_layer_0; // @[Cave.scala 166:32]
  assign gpu_io_layerCtrl_0_format = 4'h4 == gameIndexReg ? 2'h3 : _gameConfig_T_11_layer_0_format; // @[Mux.scala 81:58]
  assign gpu_io_layerCtrl_0_regs_tileSize = main_io_gpuMem_layer_0_regs_tileSize; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_0_regs_enable = main_io_gpuMem_layer_0_regs_enable; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_0_regs_flipX = main_io_gpuMem_layer_0_regs_flipX; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_0_regs_flipY = main_io_gpuMem_layer_0_regs_flipY; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_0_regs_rowScrollEnable = main_io_gpuMem_layer_0_regs_rowScrollEnable; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_0_regs_rowSelectEnable = main_io_gpuMem_layer_0_regs_rowSelectEnable; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_0_regs_scroll_x = main_io_gpuMem_layer_0_regs_scroll_x; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_0_regs_scroll_y = main_io_gpuMem_layer_0_regs_scroll_y; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_0_vram8x8_dout = main_io_gpuMem_layer_0_vram8x8_dout; // @[Cave.scala 168:33]
  assign gpu_io_layerCtrl_0_vram16x16_dout = main_io_gpuMem_layer_0_vram16x16_dout; // @[Cave.scala 169:35]
  assign gpu_io_layerCtrl_0_lineRam_dout = main_io_gpuMem_layer_0_lineRam_dout; // @[Cave.scala 170:33]
  assign gpu_io_layerCtrl_0_tileRom_dout = gpu_io_layerCtrl_0_tileRom_crossing_io_in_dout; // @[Cave.scala 171:33]
  assign gpu_io_layerCtrl_1_enable = options_layer_1; // @[Cave.scala 166:32]
  assign gpu_io_layerCtrl_1_format = 4'h4 == gameIndexReg ? 2'h0 : _gameConfig_T_11_layer_0_format; // @[Mux.scala 81:58]
  assign gpu_io_layerCtrl_1_regs_tileSize = main_io_gpuMem_layer_1_regs_tileSize; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_1_regs_enable = main_io_gpuMem_layer_1_regs_enable; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_1_regs_flipX = main_io_gpuMem_layer_1_regs_flipX; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_1_regs_flipY = main_io_gpuMem_layer_1_regs_flipY; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_1_regs_rowScrollEnable = main_io_gpuMem_layer_1_regs_rowScrollEnable; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_1_regs_rowSelectEnable = main_io_gpuMem_layer_1_regs_rowSelectEnable; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_1_regs_scroll_x = main_io_gpuMem_layer_1_regs_scroll_x; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_1_regs_scroll_y = main_io_gpuMem_layer_1_regs_scroll_y; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_1_vram8x8_dout = main_io_gpuMem_layer_1_vram8x8_dout; // @[Cave.scala 168:33]
  assign gpu_io_layerCtrl_1_vram16x16_dout = main_io_gpuMem_layer_1_vram16x16_dout; // @[Cave.scala 169:35]
  assign gpu_io_layerCtrl_1_lineRam_dout = main_io_gpuMem_layer_1_lineRam_dout; // @[Cave.scala 170:33]
  assign gpu_io_layerCtrl_1_tileRom_dout = gpu_io_layerCtrl_1_tileRom_crossing_io_in_dout; // @[Cave.scala 171:33]
  assign gpu_io_layerCtrl_2_enable = options_layer_2; // @[Cave.scala 166:32]
  assign gpu_io_layerCtrl_2_format = 4'h4 == gameIndexReg ? 2'h0 : _gameConfig_T_11_layer_2_format; // @[Mux.scala 81:58]
  assign gpu_io_layerCtrl_2_regs_tileSize = main_io_gpuMem_layer_2_regs_tileSize; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_2_regs_enable = main_io_gpuMem_layer_2_regs_enable; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_2_regs_flipX = main_io_gpuMem_layer_2_regs_flipX; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_2_regs_flipY = main_io_gpuMem_layer_2_regs_flipY; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_2_regs_rowScrollEnable = main_io_gpuMem_layer_2_regs_rowScrollEnable; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_2_regs_rowSelectEnable = main_io_gpuMem_layer_2_regs_rowSelectEnable; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_2_regs_scroll_x = main_io_gpuMem_layer_2_regs_scroll_x; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_2_regs_scroll_y = main_io_gpuMem_layer_2_regs_scroll_y; // @[Cave.scala 172:30]
  assign gpu_io_layerCtrl_2_vram8x8_dout = main_io_gpuMem_layer_2_vram8x8_dout; // @[Cave.scala 168:33]
  assign gpu_io_layerCtrl_2_vram16x16_dout = main_io_gpuMem_layer_2_vram16x16_dout; // @[Cave.scala 169:35]
  assign gpu_io_layerCtrl_2_lineRam_dout = main_io_gpuMem_layer_2_lineRam_dout; // @[Cave.scala 170:33]
  assign gpu_io_layerCtrl_2_tileRom_dout = gpu_io_layerCtrl_2_tileRom_crossing_io_in_dout; // @[Cave.scala 171:33]
  assign gpu_io_spriteCtrl_enable = options_sprite; // @[Cave.scala 174:28]
  assign gpu_io_spriteCtrl_format = 4'h4 == gameIndexReg ? 2'h1 : _gameConfig_T_11_sprite_format; // @[Mux.scala 81:58]
  assign gpu_io_spriteCtrl_start = ~vBlank & vBlankFalling_REG; // @[Util.scala 165:35]
  assign gpu_io_spriteCtrl_zoom = 4'h4 == gameIndexReg | (4'h7 == gameIndexReg | (4'h5 == gameIndexReg | (4'h6 ==
    gameIndexReg | (4'h3 == gameIndexReg | _gameConfig_T_3_sprite_zoom)))); // @[Mux.scala 81:58]
  assign gpu_io_spriteCtrl_regs_offset_x = main_io_gpuMem_sprite_regs_offset_x; // @[Cave.scala 180:26]
  assign gpu_io_spriteCtrl_regs_offset_y = main_io_gpuMem_sprite_regs_offset_y; // @[Cave.scala 180:26]
  assign gpu_io_spriteCtrl_regs_bank = main_io_gpuMem_sprite_regs_bank; // @[Cave.scala 180:26]
  assign gpu_io_spriteCtrl_regs_fixed = main_io_gpuMem_sprite_regs_fixed; // @[Cave.scala 180:26]
  assign gpu_io_spriteCtrl_regs_hFlip = main_io_gpuMem_sprite_regs_hFlip; // @[Cave.scala 180:26]
  assign gpu_io_spriteCtrl_vram_dout = main_io_gpuMem_sprite_vram_dout; // @[Cave.scala 178:26]
  assign gpu_io_spriteCtrl_tileRom_dout = memSys_io_spriteTileRom_dout; // @[Cave.scala 179:29]
  assign gpu_io_spriteCtrl_tileRom_wait_n = memSys_io_spriteTileRom_wait_n; // @[Cave.scala 179:29]
  assign gpu_io_spriteCtrl_tileRom_valid = memSys_io_spriteTileRom_valid; // @[Cave.scala 179:29]
  assign gpu_io_spriteCtrl_tileRom_burstDone = memSys_io_spriteTileRom_burstDone; // @[Cave.scala 179:29]
  assign gpu_io_gameConfig_granularity = 4'h4 == gameIndexReg ? 9'h100 : _gameConfig_T_11_granularity; // @[Mux.scala 81:58]
  assign gpu_io_gameConfig_layer_0_paletteBank = 4'h4 == gameIndexReg ? 2'h1 : _gameConfig_T_11_layer_0_paletteBank; // @[Mux.scala 81:58]
  assign gpu_io_gameConfig_layer_1_paletteBank = 4'h4 == gameIndexReg ? 2'h0 : _gameConfig_T_11_layer_0_paletteBank; // @[Mux.scala 81:58]
  assign gpu_io_gameConfig_layer_2_paletteBank = 4'h4 == gameIndexReg ? 2'h0 : _gameConfig_T_11_layer_2_paletteBank; // @[Mux.scala 81:58]
  assign gpu_io_options_rotate = options_rotate; // @[Cave.scala 182:18]
  assign gpu_io_options_flip = options_flip; // @[Cave.scala 182:18]
  assign gpu_io_video_clockEnable = videoSys_io_video_clockEnable; // @[Cave.scala 183:16]
  assign gpu_io_video_displayEnable = videoSys_io_video_displayEnable; // @[Cave.scala 183:16]
  assign gpu_io_video_pos_x = videoSys_io_video_pos_x; // @[Cave.scala 183:16]
  assign gpu_io_video_pos_y = videoSys_io_video_pos_y; // @[Cave.scala 183:16]
  assign gpu_io_video_vBlank = videoSys_io_video_vBlank; // @[Cave.scala 183:16]
  assign gpu_io_video_regs_size_x = videoSys_io_video_regs_size_x; // @[Cave.scala 183:16]
  assign gpu_io_video_regs_size_y = videoSys_io_video_regs_size_y; // @[Cave.scala 183:16]
  assign gpu_io_spriteLineBuffer_dout = spriteFrameBuffer_io_lineBuffer_dout; // @[Cave.scala 192:35]
  assign gpu_io_spriteFrameBuffer_wait_n = spriteFrameBuffer_io_frameBuffer_wait_n; // @[Cave.scala 193:36]
  assign gpu_io_paletteRam_dout = main_io_gpuMem_paletteRam_dout; // @[Cave.scala 184:21]
  assign gpu_io_layerCtrl_0_tileRom_crossing_clock = clock;
  assign gpu_io_layerCtrl_0_tileRom_crossing_io_targetClock = videoClock; // @[Crossing.scala 201:29]
  assign gpu_io_layerCtrl_0_tileRom_crossing_io_in_rd = gpu_io_layerCtrl_0_tileRom_rd; // @[Cave.scala 171:33]
  assign gpu_io_layerCtrl_0_tileRom_crossing_io_in_addr = gpu_io_layerCtrl_0_tileRom_addr; // @[Cave.scala 171:33]
  assign gpu_io_layerCtrl_0_tileRom_crossing_io_out_dout = memSys_io_layerTileRom_0_dout; // @[Crossing.scala 202:21]
  assign gpu_io_layerCtrl_0_tileRom_crossing_io_out_wait_n = memSys_io_layerTileRom_0_wait_n; // @[Crossing.scala 202:21]
  assign gpu_io_layerCtrl_0_tileRom_crossing_io_out_valid = memSys_io_layerTileRom_0_valid; // @[Crossing.scala 202:21]
  assign gpu_io_layerCtrl_1_tileRom_crossing_clock = clock;
  assign gpu_io_layerCtrl_1_tileRom_crossing_io_targetClock = videoClock; // @[Crossing.scala 201:29]
  assign gpu_io_layerCtrl_1_tileRom_crossing_io_in_rd = gpu_io_layerCtrl_1_tileRom_rd; // @[Cave.scala 171:33]
  assign gpu_io_layerCtrl_1_tileRom_crossing_io_in_addr = gpu_io_layerCtrl_1_tileRom_addr; // @[Cave.scala 171:33]
  assign gpu_io_layerCtrl_1_tileRom_crossing_io_out_dout = memSys_io_layerTileRom_1_dout; // @[Crossing.scala 202:21]
  assign gpu_io_layerCtrl_1_tileRom_crossing_io_out_wait_n = memSys_io_layerTileRom_1_wait_n; // @[Crossing.scala 202:21]
  assign gpu_io_layerCtrl_1_tileRom_crossing_io_out_valid = memSys_io_layerTileRom_1_valid; // @[Crossing.scala 202:21]
  assign gpu_io_layerCtrl_2_tileRom_crossing_clock = clock;
  assign gpu_io_layerCtrl_2_tileRom_crossing_io_targetClock = videoClock; // @[Crossing.scala 201:29]
  assign gpu_io_layerCtrl_2_tileRom_crossing_io_in_rd = gpu_io_layerCtrl_2_tileRom_rd; // @[Cave.scala 171:33]
  assign gpu_io_layerCtrl_2_tileRom_crossing_io_in_addr = gpu_io_layerCtrl_2_tileRom_addr; // @[Cave.scala 171:33]
  assign gpu_io_layerCtrl_2_tileRom_crossing_io_out_dout = memSys_io_layerTileRom_2_dout; // @[Crossing.scala 202:21]
  assign gpu_io_layerCtrl_2_tileRom_crossing_io_out_wait_n = memSys_io_layerTileRom_2_wait_n; // @[Crossing.scala 202:21]
  assign gpu_io_layerCtrl_2_tileRom_crossing_io_out_valid = memSys_io_layerTileRom_2_valid; // @[Crossing.scala 202:21]
  assign spriteFrameBuffer_clock = clock;
  assign spriteFrameBuffer_reset = reset;
  assign spriteFrameBuffer_io_videoClock = videoClock; // @[Cave.scala 188:35]
  assign spriteFrameBuffer_io_enable = memSys_io_ready; // @[Cave.scala 189:31]
  assign spriteFrameBuffer_io_swap = main_io_spriteFrameBufferSwap; // @[Cave.scala 190:29]
  assign spriteFrameBuffer_io_video_pos_y = videoSys_io_video_pos_y; // @[Cave.scala 191:30]
  assign spriteFrameBuffer_io_video_hBlank = videoSys_io_video_hBlank; // @[Cave.scala 191:30]
  assign spriteFrameBuffer_io_lineBuffer_addr = gpu_io_spriteLineBuffer_addr; // @[Cave.scala 192:35]
  assign spriteFrameBuffer_io_frameBuffer_wr = gpu_io_spriteFrameBuffer_wr; // @[Cave.scala 193:36]
  assign spriteFrameBuffer_io_frameBuffer_addr = gpu_io_spriteFrameBuffer_addr; // @[Cave.scala 193:36]
  assign spriteFrameBuffer_io_frameBuffer_din = gpu_io_spriteFrameBuffer_din; // @[Cave.scala 193:36]
  assign spriteFrameBuffer_io_ddr_dout = memSys_io_spriteFrameBuffer_dout; // @[Cave.scala 194:28]
  assign spriteFrameBuffer_io_ddr_wait_n = memSys_io_spriteFrameBuffer_wait_n; // @[Cave.scala 194:28]
  assign spriteFrameBuffer_io_ddr_valid = memSys_io_spriteFrameBuffer_valid; // @[Cave.scala 194:28]
  assign spriteFrameBuffer_io_ddr_burstDone = memSys_io_spriteFrameBuffer_burstDone; // @[Cave.scala 194:28]
  assign systemFrameBuffer_clock = clock;
  assign systemFrameBuffer_reset = reset;
  assign systemFrameBuffer_io_videoClock = videoClock; // @[Cave.scala 198:35]
  assign systemFrameBuffer_io_enable = memSys_io_ready; // @[Cave.scala 199:31]
  assign systemFrameBuffer_io_rotate = options_rotate; // @[Cave.scala 200:31]
  assign systemFrameBuffer_io_forceBlank = ~memSys_io_ready; // @[Cave.scala 201:38]
  assign systemFrameBuffer_io_video_vBlank = videoSys_io_video_vBlank; // @[Cave.scala 202:30]
  assign systemFrameBuffer_io_video_regs_size_x = videoSys_io_video_regs_size_x; // @[Cave.scala 202:30]
  assign systemFrameBuffer_io_video_regs_size_y = videoSys_io_video_regs_size_y; // @[Cave.scala 202:30]
  assign systemFrameBuffer_io_frameBufferCtrl_vBlank = frameBufferCtrl_vBlank; // @[Cave.scala 203:40]
  assign systemFrameBuffer_io_frameBufferCtrl_lowLat = frameBufferCtrl_lowLat; // @[Cave.scala 203:40]
  assign systemFrameBuffer_io_frameBuffer_wr = gpu_io_systemFrameBuffer_wr; // @[Cave.scala 204:36]
  assign systemFrameBuffer_io_frameBuffer_addr = gpu_io_systemFrameBuffer_addr; // @[Cave.scala 204:36]
  assign systemFrameBuffer_io_frameBuffer_din = gpu_io_systemFrameBuffer_din; // @[Cave.scala 204:36]
  assign systemFrameBuffer_io_ddr_wait_n = memSys_io_systemFrameBuffer_wait_n; // @[Cave.scala 205:28]
  always @(posedge clock) begin
    vBlank_r <= video_vBlank; // @[Reg.scala 19:16 20:{18,22}]
    vBlank <= vBlank_r; // @[Reg.scala 19:16 20:{18,22}]
    vBlankFalling_REG <= vBlank; // @[Util.scala 165:45]
    if (_gameIndexReg_T_4 & ~gameIndexReg_latched) begin // @[Cave.scala 101:55]
      gameIndexReg <= options_gameIndex; // @[Cave.scala 102:11]
    end else if (ioctl_download & ioctl_wr & ioctl_index == 8'h1) begin // @[Cave.scala 97:85]
      gameIndexReg <= ioctl_dout[3:0]; // @[Cave.scala 98:11]
    end
    if (reset) begin // @[Cave.scala 96:26]
      gameIndexReg_latched <= 1'h0; // @[Cave.scala 96:26]
    end else begin
      gameIndexReg_latched <= _GEN_5;
    end
    gameIndexReg_REG <= ioctl_download; // @[Util.scala 165:45]
    if (memSys_io_prog_nvram_mem_valid) begin // @[Reg.scala 20:18]
      memSys_io_prog_nvram_view__ioctl_din_r <= memSys_io_prog_nvram_mem_dout; // @[Reg.scala 20:22]
    end
    memSys_io_prog_done_REG <= ioctl_download; // @[Util.scala 165:45]
    videoSys_io_prog_done_REG <= ioctl_download; // @[Util.scala 165:45]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  vBlank_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  vBlank = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  vBlankFalling_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  gameIndexReg = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  gameIndexReg_latched = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  gameIndexReg_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  memSys_io_prog_nvram_view__ioctl_din_r = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  memSys_io_prog_done_REG = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  videoSys_io_prog_done_REG = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
