module SystemFrameBuffer(
  input         clock,
  input         reset,
  input         io_videoClock,
  input         io_enable,
  input         io_rotate,
  input         io_forceBlank,
  input         io_video_vBlank,
  input  [8:0]  io_video_regs_size_x,
  input  [8:0]  io_video_regs_size_y,
  output        io_frameBufferCtrl_enable,
  output [11:0] io_frameBufferCtrl_hSize,
  output [11:0] io_frameBufferCtrl_vSize,
  output [31:0] io_frameBufferCtrl_baseAddr,
  output [13:0] io_frameBufferCtrl_stride,
  input         io_frameBufferCtrl_vBlank,
  input         io_frameBufferCtrl_lowLat,
  output        io_frameBufferCtrl_forceBlank,
  input         io_frameBuffer_wr,
  input  [16:0] io_frameBuffer_addr,
  input  [31:0] io_frameBuffer_din,
  output        io_ddr_wr,
  output [31:0] io_ddr_addr,
  output [7:0]  io_ddr_mask,
  output [63:0] io_ddr_din,
  input         io_ddr_wait_n
);

  wire [31:0] _queue_io_out_addr;
  wire        _pageFlipper_io_mode;
  wire        _pageFlipper_io_swapRead;
  wire        _pageFlipper_io_swapWrite;
  wire [31:0] _pageFlipper_io_addrWrite;
  reg         pageFlipper_io_swapRead_r;
  reg         pageFlipper_io_swapRead_r_1;
  reg         pageFlipper_io_swapRead_REG;
  reg         pageFlipper_io_swapWrite_r;
  reg         pageFlipper_io_swapWrite_r_1;
  reg         pageFlipper_io_swapWrite_REG;
  wire [8:0]  _io_frameBufferCtrl_hSize_T =
    io_rotate ? io_video_regs_size_y : io_video_regs_size_x;
  wire [8:0]  _io_frameBufferCtrl_vSize_T =
    io_rotate ? io_video_regs_size_x : io_video_regs_size_y;
  wire [8:0]  _GEN = io_rotate ? io_video_regs_size_y : io_video_regs_size_x;
  always @(posedge clock) begin
    pageFlipper_io_swapRead_r <= io_frameBufferCtrl_vBlank;
    pageFlipper_io_swapRead_r_1 <= pageFlipper_io_swapRead_r;
    pageFlipper_io_swapRead_REG <= pageFlipper_io_swapRead_r_1;
    pageFlipper_io_swapWrite_r <= io_video_vBlank;
    pageFlipper_io_swapWrite_r_1 <= pageFlipper_io_swapWrite_r;
    pageFlipper_io_swapWrite_REG <= pageFlipper_io_swapWrite_r_1;
  end // always @(posedge)
  assign _pageFlipper_io_mode = ~io_frameBufferCtrl_lowLat;
  assign _pageFlipper_io_swapRead =
    pageFlipper_io_swapRead_r_1 & ~pageFlipper_io_swapRead_REG;
  assign _pageFlipper_io_swapWrite =
    pageFlipper_io_swapWrite_r_1 & ~pageFlipper_io_swapWrite_REG;
  PageFlipper_1 pageFlipper (
    .clock        (clock),
    .reset        (reset),
    .io_mode      (_pageFlipper_io_mode),
    .io_swapRead  (_pageFlipper_io_swapRead),
    .io_swapWrite (_pageFlipper_io_swapWrite),
    .io_addrRead  (io_frameBufferCtrl_baseAddr),
    .io_addrWrite (_pageFlipper_io_addrWrite)
  );
  RequestQueue_1 queue (
    .clock         (io_videoClock),
    .io_enable     (io_enable),
    .io_readClock  (clock),
    .io_in_wr      (io_frameBuffer_wr),
    .io_in_addr    (io_frameBuffer_addr),
    .io_in_din     (io_frameBuffer_din),
    .io_out_wr     (io_ddr_wr),
    .io_out_addr   (_queue_io_out_addr),
    .io_out_mask   (io_ddr_mask),
    .io_out_din    (io_ddr_din),
    .io_out_wait_n (io_ddr_wait_n)
  );
  assign io_frameBufferCtrl_enable = io_enable;
  assign io_frameBufferCtrl_hSize = {3'h0, _io_frameBufferCtrl_hSize_T};
  assign io_frameBufferCtrl_vSize = {3'h0, _io_frameBufferCtrl_vSize_T};
  assign io_frameBufferCtrl_stride = {3'h0, _GEN, 2'h0};
  assign io_frameBufferCtrl_forceBlank = io_forceBlank;
  assign io_ddr_addr = 32'(_queue_io_out_addr + _pageFlipper_io_addrWrite);
endmodule

