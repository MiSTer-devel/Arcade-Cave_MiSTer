module LayerProcessor_1(
  input         clock,
  input         io_ctrl_enable,
  input  [1:0]  io_ctrl_format,
  input         io_ctrl_regs_tileSize,
  input         io_ctrl_regs_enable,
  input         io_ctrl_regs_flipX,
  input         io_ctrl_regs_flipY,
  input         io_ctrl_regs_rowScrollEnable,
  input         io_ctrl_regs_rowSelectEnable,
  input  [8:0]  io_ctrl_regs_scroll_x,
  input  [8:0]  io_ctrl_regs_scroll_y,
  output [11:0] io_ctrl_vram8x8_addr,
  input  [31:0] io_ctrl_vram8x8_dout,
  output [9:0]  io_ctrl_vram16x16_addr,
  input  [31:0] io_ctrl_vram16x16_dout,
  output [8:0]  io_ctrl_lineRam_addr,
  input  [31:0] io_ctrl_lineRam_dout,
  output        io_ctrl_tileRom_rd,
  output [31:0] io_ctrl_tileRom_addr,
  input  [63:0] io_ctrl_tileRom_dout,
  input         io_video_clockEnable,
  input  [8:0]  io_video_pos_x,
  input  [8:0]  io_video_pos_y,
  input         io_video_vBlank,
  input  [8:0]  io_video_regs_size_x,
  input  [8:0]  io_video_regs_size_y,
  input  [8:0]  io_spriteOffset_x,
  input  [8:0]  io_spriteOffset_y,
  output [1:0]  io_pen_priority,
  output [5:0]  io_pen_palette,
  output [7:0]  io_pen_color
);

  reg  [8:0]  lineEffectReg_rowSelect;
  reg  [8:0]  lineEffectReg_rowScroll;
  wire        layerEnable = io_ctrl_enable & (|io_ctrl_format) & io_ctrl_regs_enable;
  wire [4:0]  layerOffset_x = io_ctrl_regs_tileSize ? 5'h11 : 5'h9;
  wire [4:0]  _layerOffset_T_2 =
    io_ctrl_regs_flipX ? 5'(layerOffset_x + 5'h1) : layerOffset_x;
  wire [8:0]  _GEN = {4'h0, _layerOffset_T_2};
  wire [8:0]  _GEN_0 = {8'hF7, io_ctrl_regs_flipY};
  wire [8:0]  pos_x =
    io_ctrl_regs_flipX
      ? 9'(_GEN
           + 9'(9'(9'(io_video_regs_size_x - io_video_pos_x) + io_ctrl_regs_scroll_x)
                - io_spriteOffset_x))
      : 9'(9'(9'(io_video_pos_x + io_ctrl_regs_scroll_x) - io_spriteOffset_x) - _GEN);
  wire [8:0]  pos_y =
    io_ctrl_regs_flipY
      ? 9'(9'(9'(9'(io_video_regs_size_y - io_video_pos_y) + io_ctrl_regs_scroll_y)
              - io_spriteOffset_y) + _GEN_0)
      : 9'(9'(9'(io_video_pos_y + io_ctrl_regs_scroll_y) - io_spriteOffset_y) - _GEN_0);
  wire [8:0]  _pos__x_T = io_ctrl_regs_rowScrollEnable ? lineEffectReg_rowScroll : 9'h0;
  wire [8:0]  _pos__x_T_1 = 9'(_pos__x_T + pos_x);
  wire [8:0]  pos__y = io_ctrl_regs_rowSelectEnable ? lineEffectReg_rowSelect : pos_y;
  wire [3:0]  tileOffset_x =
    io_ctrl_regs_tileSize ? _pos__x_T_1[3:0] : {1'h0, _pos__x_T_1[2:0]};
  wire [3:0]  tileOffset_y = io_ctrl_regs_tileSize ? pos__y[3:0] : {1'h0, pos__y[2:0]};
  wire [4:0]  _vramAddr_large_T_2 = io_ctrl_regs_flipX ? 5'h1F : 5'h1;
  wire [5:0]  _vramAddr_small_T_2 = io_ctrl_regs_flipX ? 6'h3F : 6'h1;
  wire [11:0] vramAddr =
    io_ctrl_regs_tileSize
      ? {2'h0, pos__y[8:4], 5'(_pos__x_T_1[8:4] + _vramAddr_large_T_2)}
      : {pos__y[8:3], 6'(_pos__x_T_1[8:3] + _vramAddr_small_T_2)};
  reg  [1:0]  tileReg_priority;
  reg  [5:0]  tileReg_colorCode;
  reg  [17:0] tileReg_code;
  reg  [1:0]  priorityReg;
  reg  [5:0]  colorReg;
  reg  [7:0]  pixReg_0;
  reg  [7:0]  pixReg_1;
  reg  [7:0]  pixReg_2;
  reg  [7:0]  pixReg_3;
  reg  [7:0]  pixReg_4;
  reg  [7:0]  pixReg_5;
  reg  [7:0]  pixReg_6;
  reg  [7:0]  pixReg_7;
  reg  [7:0]  casez_tmp;
  always @(*) begin
    casez (tileOffset_x[2:0])
      3'b000:
        casez_tmp = pixReg_0;
      3'b001:
        casez_tmp = pixReg_1;
      3'b010:
        casez_tmp = pixReg_2;
      3'b011:
        casez_tmp = pixReg_3;
      3'b100:
        casez_tmp = pixReg_4;
      3'b101:
        casez_tmp = pixReg_5;
      3'b110:
        casez_tmp = pixReg_6;
      default:
        casez_tmp = pixReg_7;
    endcase
  end // always @(*)
  wire        _io_ctrl_tileRom_addr_format16x16x4_T = io_ctrl_format == 2'h1;
  wire [25:0] _io_ctrl_tileRom_addr_T_22 =
    io_ctrl_regs_tileSize & (&io_ctrl_format)
      ? {tileReg_code, tileOffset_y[3], ~(tileOffset_x[3]), tileOffset_y[2:0], 3'h0}
      : 26'h0;
  wire [25:0] _io_ctrl_tileRom_addr_T_23 =
    io_ctrl_regs_tileSize & _io_ctrl_tileRom_addr_format16x16x4_T
      ? {1'h0, tileReg_code, tileOffset_y[3], ~(tileOffset_x[3]), tileOffset_y[2:1], 3'h0}
      : _io_ctrl_tileRom_addr_T_22;
  wire [25:0] _io_ctrl_tileRom_addr_T_24 =
    ~io_ctrl_regs_tileSize & (&io_ctrl_format)
      ? {2'h0, tileReg_code, tileOffset_y[2:0], 3'h0}
      : _io_ctrl_tileRom_addr_T_23;
  wire [25:0] _io_ctrl_tileRom_addr_T_25 =
    ~io_ctrl_regs_tileSize & _io_ctrl_tileRom_addr_format16x16x4_T
      ? {3'h0, tileReg_code, tileOffset_y[2:1], 3'h0}
      : _io_ctrl_tileRom_addr_T_24;
  wire [31:0] pixReg_pixels_4BPP_bits =
    tileOffset_y[0] ? io_ctrl_tileRom_dout[31:0] : io_ctrl_tileRom_dout[63:32];
  wire        _latchTile_T_3 =
    io_ctrl_regs_tileSize ? tileOffset_x == 4'hA : tileOffset_x == 4'h2;
  wire        _latchTile_T_4 = io_ctrl_regs_flipX ? tileOffset_x == 4'h5 : _latchTile_T_3;
  wire        _latchColor_T_3 =
    io_ctrl_regs_tileSize ? (&tileOffset_x) : tileOffset_x == 4'h7;
  wire        _latchColor_T_4 =
    io_ctrl_regs_flipX ? tileOffset_x == 4'h0 : _latchColor_T_3;
  wire        _latchPix_T_4 =
    io_ctrl_regs_flipX ? tileOffset_x[2:0] == 3'h0 : (&(tileOffset_x[2:0]));
  always @(posedge clock) begin
    if (io_video_clockEnable) begin
      lineEffectReg_rowSelect <= io_ctrl_lineRam_dout[24:16];
      lineEffectReg_rowScroll <= io_ctrl_lineRam_dout[8:0];
    end
    if (io_video_clockEnable & _latchTile_T_4) begin
      tileReg_priority <=
        io_ctrl_regs_tileSize
          ? io_ctrl_vram16x16_dout[15:14]
          : io_ctrl_vram8x8_dout[15:14];
      tileReg_colorCode <=
        io_ctrl_regs_tileSize ? io_ctrl_vram16x16_dout[13:8] : io_ctrl_vram8x8_dout[13:8];
      tileReg_code <=
        io_ctrl_regs_tileSize
          ? {2'h0, io_ctrl_vram16x16_dout[31:16]}
          : {io_ctrl_vram8x8_dout[1:0], io_ctrl_vram8x8_dout[31:16]};
    end
    if (io_video_clockEnable & _latchColor_T_4) begin
      priorityReg <= tileReg_priority;
      colorReg <= tileReg_colorCode;
    end
    if (io_video_clockEnable & _latchPix_T_4) begin
      pixReg_0 <=
        (&io_ctrl_format)
          ? {io_ctrl_tileRom_dout[55:52], io_ctrl_tileRom_dout[63:60]}
          : {4'h0, pixReg_pixels_4BPP_bits[31:28]};
      pixReg_1 <=
        (&io_ctrl_format)
          ? {io_ctrl_tileRom_dout[51:48], io_ctrl_tileRom_dout[59:56]}
          : {4'h0, pixReg_pixels_4BPP_bits[27:24]};
      pixReg_2 <=
        (&io_ctrl_format)
          ? {io_ctrl_tileRom_dout[39:36], io_ctrl_tileRom_dout[47:44]}
          : {4'h0, pixReg_pixels_4BPP_bits[23:20]};
      pixReg_3 <=
        (&io_ctrl_format)
          ? {io_ctrl_tileRom_dout[35:32], io_ctrl_tileRom_dout[43:40]}
          : {4'h0, pixReg_pixels_4BPP_bits[19:16]};
      pixReg_4 <=
        (&io_ctrl_format)
          ? {io_ctrl_tileRom_dout[23:20], io_ctrl_tileRom_dout[31:28]}
          : {4'h0, pixReg_pixels_4BPP_bits[15:12]};
      pixReg_5 <=
        (&io_ctrl_format)
          ? {io_ctrl_tileRom_dout[19:16], io_ctrl_tileRom_dout[27:24]}
          : {4'h0, pixReg_pixels_4BPP_bits[11:8]};
      pixReg_6 <=
        (&io_ctrl_format)
          ? {io_ctrl_tileRom_dout[7:4], io_ctrl_tileRom_dout[15:12]}
          : {4'h0, pixReg_pixels_4BPP_bits[7:4]};
      pixReg_7 <=
        (&io_ctrl_format)
          ? {io_ctrl_tileRom_dout[3:0], io_ctrl_tileRom_dout[11:8]}
          : {4'h0, pixReg_pixels_4BPP_bits[3:0]};
    end
  end // always @(posedge)
  assign io_ctrl_vram8x8_addr = vramAddr;
  assign io_ctrl_vram16x16_addr = vramAddr[9:0];
  assign io_ctrl_lineRam_addr = io_ctrl_regs_flipY ? 9'(pos_y + 9'h1) : 9'(pos_y - 9'h1);
  assign io_ctrl_tileRom_rd = layerEnable & ~io_video_vBlank;
  assign io_ctrl_tileRom_addr = {6'h0, _io_ctrl_tileRom_addr_T_25};
  assign io_pen_priority = layerEnable ? priorityReg : 2'h0;
  assign io_pen_palette = layerEnable ? colorReg : 6'h0;
  assign io_pen_color = layerEnable ? casez_tmp : 8'h0;
endmodule

