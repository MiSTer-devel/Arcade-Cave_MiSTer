module MemSys(
  input         clock,
  input         reset,
  input  [31:0] io_gameConfig_eepromOffset,
  input  [31:0] io_gameConfig_sound_0_romOffset,
  input  [31:0] io_gameConfig_sound_1_romOffset,
  input  [31:0] io_gameConfig_layer_0_romOffset,
  input  [31:0] io_gameConfig_layer_1_romOffset,
  input  [31:0] io_gameConfig_layer_2_romOffset,
  input  [31:0] io_gameConfig_sprite_romOffset,
  input         io_prog_rom_wr,
  input  [26:0] io_prog_rom_addr,
  input  [15:0] io_prog_rom_din,
  output        io_prog_rom_wait_n,
  input         io_prog_nvram_rd,
  input         io_prog_nvram_wr,
  input  [26:0] io_prog_nvram_addr,
  input  [15:0] io_prog_nvram_din,
  output [15:0] io_prog_nvram_dout,
  output        io_prog_nvram_wait_n,
  output        io_prog_nvram_valid,
  input         io_prog_done,
  input         io_progRom_rd,
  input  [19:0] io_progRom_addr,
  output [15:0] io_progRom_dout,
  output        io_progRom_wait_n,
  output        io_progRom_valid,
  input         io_eeprom_rd,
  input         io_eeprom_wr,
  input  [6:0]  io_eeprom_addr,
  input  [15:0] io_eeprom_din,
  output [15:0] io_eeprom_dout,
  output        io_eeprom_wait_n,
  output        io_eeprom_valid,
  input         io_soundRom_0_rd,
  input  [24:0] io_soundRom_0_addr,
  output [7:0]  io_soundRom_0_dout,
  output        io_soundRom_0_wait_n,
  output        io_soundRom_0_valid,
  input         io_soundRom_1_rd,
  input  [24:0] io_soundRom_1_addr,
  output [7:0]  io_soundRom_1_dout,
  output        io_soundRom_1_wait_n,
  output        io_soundRom_1_valid,
  input         io_layerTileRom_0_rd,
  input  [31:0] io_layerTileRom_0_addr,
  output [63:0] io_layerTileRom_0_dout,
  output        io_layerTileRom_0_wait_n,
  output        io_layerTileRom_0_valid,
  input         io_layerTileRom_1_rd,
  input  [31:0] io_layerTileRom_1_addr,
  output [63:0] io_layerTileRom_1_dout,
  output        io_layerTileRom_1_wait_n,
  output        io_layerTileRom_1_valid,
  input         io_layerTileRom_2_rd,
  input  [31:0] io_layerTileRom_2_addr,
  output [63:0] io_layerTileRom_2_dout,
  output        io_layerTileRom_2_wait_n,
  output        io_layerTileRom_2_valid,
  input         io_spriteTileRom_rd,
  input  [31:0] io_spriteTileRom_addr,
  output [63:0] io_spriteTileRom_dout,
  output        io_spriteTileRom_wait_n,
  output        io_spriteTileRom_valid,
  input  [7:0]  io_spriteTileRom_burstLength,
  output        io_spriteTileRom_burstDone,
  output        io_ddr_rd,
  output        io_ddr_wr,
  output [31:0] io_ddr_addr,
  output [7:0]  io_ddr_mask,
  output [63:0] io_ddr_din,
  input  [63:0] io_ddr_dout,
  input         io_ddr_wait_n,
  input         io_ddr_valid,
  output [7:0]  io_ddr_burstLength,
  input         io_ddr_burstDone,
  output        io_sdram_rd,
  output        io_sdram_wr,
  output [24:0] io_sdram_addr,
  output [15:0] io_sdram_din,
  input  [15:0] io_sdram_dout,
  input         io_sdram_wait_n,
  input         io_sdram_valid,
  input         io_sdram_burstDone,
  input         io_spriteFrameBuffer_rd,
  input         io_spriteFrameBuffer_wr,
  input  [31:0] io_spriteFrameBuffer_addr,
  input  [7:0]  io_spriteFrameBuffer_mask,
  input  [63:0] io_spriteFrameBuffer_din,
  output [63:0] io_spriteFrameBuffer_dout,
  output        io_spriteFrameBuffer_wait_n,
  output        io_spriteFrameBuffer_valid,
  input  [7:0]  io_spriteFrameBuffer_burstLength,
  output        io_spriteFrameBuffer_burstDone,
  input         io_systemFrameBuffer_wr,
  input  [31:0] io_systemFrameBuffer_addr,
  input  [7:0]  io_systemFrameBuffer_mask,
  input  [63:0] io_systemFrameBuffer_din,
  output        io_systemFrameBuffer_wait_n,
  output        io_ready
);

  reg         io_ready_enableReg;
  wire [6:0]  _nvramArbiter_io_in_0_addr;
  wire [24:0] _sdramArbiter_io_in_2_addr;
  wire [24:0] _sdramArbiter_io_in_3_addr;
  wire [24:0] _sdramArbiter_io_in_4_addr;
  wire [24:0] _sdramArbiter_io_in_5_addr;
  wire [24:0] _sdramArbiter_io_in_6_addr;
  wire [24:0] _sdramArbiter_io_in_7_addr;
  wire [31:0] _ddrArbiter_io_in_0_addr;
  wire [31:0] _ddrArbiter_io_in_1_addr;
  wire [31:0] _ddrArbiter_io_in_4_addr;
  wire [15:0] _layerRomCache_2_io_out_dout;
  wire        _layerRomCache_2_io_out_wait_n;
  wire        _layerRomCache_2_io_out_valid;
  wire        _layerRomCache_2_io_out_rd;
  wire [24:0] _layerRomCache_2_io_out_addr;
  wire [15:0] _layerRomCache_1_io_out_dout;
  wire        _layerRomCache_1_io_out_wait_n;
  wire        _layerRomCache_1_io_out_valid;
  wire        _layerRomCache_1_io_out_rd;
  wire [24:0] _layerRomCache_1_io_out_addr;
  wire [15:0] _layerRomCache_0_io_out_dout;
  wire        _layerRomCache_0_io_out_wait_n;
  wire        _layerRomCache_0_io_out_valid;
  wire        _layerRomCache_0_io_out_rd;
  wire [24:0] _layerRomCache_0_io_out_addr;
  wire [15:0] _soundRomCache_1_io_out_dout;
  wire        _soundRomCache_1_io_out_wait_n;
  wire        _soundRomCache_1_io_out_valid;
  wire        _soundRomCache_1_io_out_rd;
  wire [24:0] _soundRomCache_1_io_out_addr;
  wire [15:0] _soundRomCache_0_io_out_dout;
  wire        _soundRomCache_0_io_out_wait_n;
  wire        _soundRomCache_0_io_out_valid;
  wire        _soundRomCache_0_io_out_rd;
  wire [24:0] _soundRomCache_0_io_out_addr;
  wire        _eepromCache_io_in_rd;
  wire        _eepromCache_io_in_wr;
  wire [6:0]  _eepromCache_io_in_addr;
  wire [15:0] _eepromCache_io_in_din;
  wire [15:0] _eepromCache_io_out_dout;
  wire        _eepromCache_io_out_wait_n;
  wire        _eepromCache_io_out_valid;
  wire [15:0] _eepromCache_io_in_dout;
  wire        _eepromCache_io_in_wait_n;
  wire        _eepromCache_io_in_valid;
  wire        _eepromCache_io_out_rd;
  wire        _eepromCache_io_out_wr;
  wire [24:0] _eepromCache_io_out_addr;
  wire [15:0] _eepromCache_io_out_din;
  wire [15:0] _progRomCache_io_out_dout;
  wire        _progRomCache_io_out_wait_n;
  wire        _progRomCache_io_out_valid;
  wire        _progRomCache_io_out_rd;
  wire [24:0] _progRomCache_io_out_addr;
  wire        _copyDma_io_start;
  wire [63:0] _copyDma_io_in_dout;
  wire        _copyDma_io_in_wait_n;
  wire        _copyDma_io_in_valid;
  wire        _copyDma_io_in_burstDone;
  wire        _copyDma_io_busy;
  wire        _copyDma_io_in_rd;
  wire [31:0] _copyDma_io_in_addr;
  wire        _sdramDownloadBuffer_io_in_wr;
  wire [31:0] _sdramDownloadBuffer_io_in_addr;
  wire [63:0] _sdramDownloadBuffer_io_in_din;
  wire        _sdramDownloadBuffer_io_out_wait_n;
  wire        _sdramDownloadBuffer_io_out_burstDone;
  wire        _sdramDownloadBuffer_io_in_wait_n;
  wire        _sdramDownloadBuffer_io_out_wr;
  wire [24:0] _sdramDownloadBuffer_io_out_addr;
  wire [15:0] _sdramDownloadBuffer_io_out_din;
  wire        _ddrDownloadBuffer_io_out_burstDone;
  wire        _ddrDownloadBuffer_io_out_wr;
  wire [31:0] _ddrDownloadBuffer_io_out_addr;
  wire [63:0] _ddrDownloadBuffer_io_out_din;
  reg         io_ready_REG;
  always @(posedge clock) begin
    io_ready_REG <= _copyDma_io_busy;
    if (reset)
      io_ready_enableReg <= 1'h0;
    else
      io_ready_enableReg <= ~_copyDma_io_busy & io_ready_REG | io_ready_enableReg;
  end // always @(posedge)
  BurstBuffer ddrDownloadBuffer (
    .clock            (clock),
    .reset            (reset),
    .io_in_wr         (io_prog_rom_wr),
    .io_in_addr       (io_prog_rom_addr),
    .io_in_din        (io_prog_rom_din),
    .io_out_wr        (_ddrDownloadBuffer_io_out_wr),
    .io_out_addr      (_ddrDownloadBuffer_io_out_addr),
    .io_out_din       (_ddrDownloadBuffer_io_out_din),
    .io_out_burstDone (_ddrDownloadBuffer_io_out_burstDone)
  );
  BurstBuffer_1 sdramDownloadBuffer (
    .clock            (clock),
    .reset            (reset),
    .io_in_wr         (_sdramDownloadBuffer_io_in_wr),
    .io_in_addr       (_sdramDownloadBuffer_io_in_addr),
    .io_in_din        (_sdramDownloadBuffer_io_in_din),
    .io_in_wait_n     (_sdramDownloadBuffer_io_in_wait_n),
    .io_out_wr        (_sdramDownloadBuffer_io_out_wr),
    .io_out_addr      (_sdramDownloadBuffer_io_out_addr),
    .io_out_din       (_sdramDownloadBuffer_io_out_din),
    .io_out_wait_n    (_sdramDownloadBuffer_io_out_wait_n),
    .io_out_burstDone (_sdramDownloadBuffer_io_out_burstDone)
  );
  assign _copyDma_io_start = ~io_ready_enableReg & io_prog_done;
  BurstReadDMA copyDma (
    .clock           (clock),
    .reset           (reset),
    .io_start        (_copyDma_io_start),
    .io_busy         (_copyDma_io_busy),
    .io_in_rd        (_copyDma_io_in_rd),
    .io_in_addr      (_copyDma_io_in_addr),
    .io_in_dout      (_copyDma_io_in_dout),
    .io_in_wait_n    (_copyDma_io_in_wait_n),
    .io_in_valid     (_copyDma_io_in_valid),
    .io_in_burstDone (_copyDma_io_in_burstDone),
    .io_out_wr       (_sdramDownloadBuffer_io_in_wr),
    .io_out_addr     (_sdramDownloadBuffer_io_in_addr),
    .io_out_din      (_sdramDownloadBuffer_io_in_din),
    .io_out_wait_n   (_sdramDownloadBuffer_io_in_wait_n)
  );
  ReadCache progRomCache (
    .clock         (clock),
    .reset         (reset),
    .io_enable     (io_ready_enableReg),
    .io_in_rd      (io_progRom_rd),
    .io_in_addr    (io_progRom_addr),
    .io_in_dout    (io_progRom_dout),
    .io_in_wait_n  (io_progRom_wait_n),
    .io_in_valid   (io_progRom_valid),
    .io_out_rd     (_progRomCache_io_out_rd),
    .io_out_addr   (_progRomCache_io_out_addr),
    .io_out_dout   (_progRomCache_io_out_dout),
    .io_out_wait_n (_progRomCache_io_out_wait_n),
    .io_out_valid  (_progRomCache_io_out_valid)
  );
  Cache eepromCache (
    .clock         (clock),
    .reset         (reset),
    .io_enable     (io_ready_enableReg),
    .io_in_rd      (_eepromCache_io_in_rd),
    .io_in_wr      (_eepromCache_io_in_wr),
    .io_in_addr    (_eepromCache_io_in_addr),
    .io_in_din     (_eepromCache_io_in_din),
    .io_in_dout    (_eepromCache_io_in_dout),
    .io_in_wait_n  (_eepromCache_io_in_wait_n),
    .io_in_valid   (_eepromCache_io_in_valid),
    .io_out_rd     (_eepromCache_io_out_rd),
    .io_out_wr     (_eepromCache_io_out_wr),
    .io_out_addr   (_eepromCache_io_out_addr),
    .io_out_din    (_eepromCache_io_out_din),
    .io_out_dout   (_eepromCache_io_out_dout),
    .io_out_wait_n (_eepromCache_io_out_wait_n),
    .io_out_valid  (_eepromCache_io_out_valid)
  );
  ReadCache_1 soundRomCache_0 (
    .clock         (clock),
    .reset         (reset),
    .io_enable     (io_ready_enableReg),
    .io_in_rd      (io_soundRom_0_rd),
    .io_in_addr    (io_soundRom_0_addr),
    .io_in_dout    (io_soundRom_0_dout),
    .io_in_wait_n  (io_soundRom_0_wait_n),
    .io_in_valid   (io_soundRom_0_valid),
    .io_out_rd     (_soundRomCache_0_io_out_rd),
    .io_out_addr   (_soundRomCache_0_io_out_addr),
    .io_out_dout   (_soundRomCache_0_io_out_dout),
    .io_out_wait_n (_soundRomCache_0_io_out_wait_n),
    .io_out_valid  (_soundRomCache_0_io_out_valid)
  );
  ReadCache_1 soundRomCache_1 (
    .clock         (clock),
    .reset         (reset),
    .io_enable     (io_ready_enableReg),
    .io_in_rd      (io_soundRom_1_rd),
    .io_in_addr    (io_soundRom_1_addr),
    .io_in_dout    (io_soundRom_1_dout),
    .io_in_wait_n  (io_soundRom_1_wait_n),
    .io_in_valid   (io_soundRom_1_valid),
    .io_out_rd     (_soundRomCache_1_io_out_rd),
    .io_out_addr   (_soundRomCache_1_io_out_addr),
    .io_out_dout   (_soundRomCache_1_io_out_dout),
    .io_out_wait_n (_soundRomCache_1_io_out_wait_n),
    .io_out_valid  (_soundRomCache_1_io_out_valid)
  );
  ReadCache_3 layerRomCache_0 (
    .clock         (clock),
    .reset         (reset),
    .io_enable     (io_ready_enableReg),
    .io_in_rd      (io_layerTileRom_0_rd),
    .io_in_addr    (io_layerTileRom_0_addr),
    .io_in_dout    (io_layerTileRom_0_dout),
    .io_in_wait_n  (io_layerTileRom_0_wait_n),
    .io_in_valid   (io_layerTileRom_0_valid),
    .io_out_rd     (_layerRomCache_0_io_out_rd),
    .io_out_addr   (_layerRomCache_0_io_out_addr),
    .io_out_dout   (_layerRomCache_0_io_out_dout),
    .io_out_wait_n (_layerRomCache_0_io_out_wait_n),
    .io_out_valid  (_layerRomCache_0_io_out_valid)
  );
  ReadCache_3 layerRomCache_1 (
    .clock         (clock),
    .reset         (reset),
    .io_enable     (io_ready_enableReg),
    .io_in_rd      (io_layerTileRom_1_rd),
    .io_in_addr    (io_layerTileRom_1_addr),
    .io_in_dout    (io_layerTileRom_1_dout),
    .io_in_wait_n  (io_layerTileRom_1_wait_n),
    .io_in_valid   (io_layerTileRom_1_valid),
    .io_out_rd     (_layerRomCache_1_io_out_rd),
    .io_out_addr   (_layerRomCache_1_io_out_addr),
    .io_out_dout   (_layerRomCache_1_io_out_dout),
    .io_out_wait_n (_layerRomCache_1_io_out_wait_n),
    .io_out_valid  (_layerRomCache_1_io_out_valid)
  );
  ReadCache_3 layerRomCache_2 (
    .clock         (clock),
    .reset         (reset),
    .io_enable     (io_ready_enableReg),
    .io_in_rd      (io_layerTileRom_2_rd),
    .io_in_addr    (io_layerTileRom_2_addr),
    .io_in_dout    (io_layerTileRom_2_dout),
    .io_in_wait_n  (io_layerTileRom_2_wait_n),
    .io_in_valid   (io_layerTileRom_2_valid),
    .io_out_rd     (_layerRomCache_2_io_out_rd),
    .io_out_addr   (_layerRomCache_2_io_out_addr),
    .io_out_dout   (_layerRomCache_2_io_out_dout),
    .io_out_wait_n (_layerRomCache_2_io_out_wait_n),
    .io_out_valid  (_layerRomCache_2_io_out_valid)
  );
  assign _ddrArbiter_io_in_0_addr = 32'(_ddrDownloadBuffer_io_out_addr + 32'h30000000);
  assign _ddrArbiter_io_in_1_addr = 32'(_copyDma_io_in_addr + 32'h30000000);
  assign _ddrArbiter_io_in_4_addr =
    32'(io_spriteTileRom_addr + 32'(io_gameConfig_sprite_romOffset + 32'h30000000));
  BurstMemArbiter ddrArbiter (
    .clock               (clock),
    .reset               (reset),
    .io_in_0_wr          (_ddrDownloadBuffer_io_out_wr),
    .io_in_0_addr        (_ddrArbiter_io_in_0_addr),
    .io_in_0_din         (_ddrDownloadBuffer_io_out_din),
    .io_in_0_burstDone   (_ddrDownloadBuffer_io_out_burstDone),
    .io_in_1_rd          (_copyDma_io_in_rd),
    .io_in_1_addr        (_ddrArbiter_io_in_1_addr),
    .io_in_1_dout        (_copyDma_io_in_dout),
    .io_in_1_wait_n      (_copyDma_io_in_wait_n),
    .io_in_1_valid       (_copyDma_io_in_valid),
    .io_in_1_burstDone   (_copyDma_io_in_burstDone),
    .io_in_2_wr          (io_systemFrameBuffer_wr),
    .io_in_2_addr        (io_systemFrameBuffer_addr),
    .io_in_2_mask        (io_systemFrameBuffer_mask),
    .io_in_2_din         (io_systemFrameBuffer_din),
    .io_in_2_wait_n      (io_systemFrameBuffer_wait_n),
    .io_in_3_rd          (io_spriteFrameBuffer_rd),
    .io_in_3_wr          (io_spriteFrameBuffer_wr),
    .io_in_3_addr        (io_spriteFrameBuffer_addr),
    .io_in_3_mask        (io_spriteFrameBuffer_mask),
    .io_in_3_din         (io_spriteFrameBuffer_din),
    .io_in_3_dout        (io_spriteFrameBuffer_dout),
    .io_in_3_wait_n      (io_spriteFrameBuffer_wait_n),
    .io_in_3_valid       (io_spriteFrameBuffer_valid),
    .io_in_3_burstLength (io_spriteFrameBuffer_burstLength),
    .io_in_3_burstDone   (io_spriteFrameBuffer_burstDone),
    .io_in_4_rd          (io_spriteTileRom_rd),
    .io_in_4_addr        (_ddrArbiter_io_in_4_addr),
    .io_in_4_dout        (io_spriteTileRom_dout),
    .io_in_4_wait_n      (io_spriteTileRom_wait_n),
    .io_in_4_valid       (io_spriteTileRom_valid),
    .io_in_4_burstLength (io_spriteTileRom_burstLength),
    .io_in_4_burstDone   (io_spriteTileRom_burstDone),
    .io_out_rd           (io_ddr_rd),
    .io_out_wr           (io_ddr_wr),
    .io_out_addr         (io_ddr_addr),
    .io_out_mask         (io_ddr_mask),
    .io_out_din          (io_ddr_din),
    .io_out_dout         (io_ddr_dout),
    .io_out_wait_n       (io_ddr_wait_n),
    .io_out_valid        (io_ddr_valid),
    .io_out_burstLength  (io_ddr_burstLength),
    .io_out_burstDone    (io_ddr_burstDone)
  );
  assign _sdramArbiter_io_in_2_addr =
    25'(_eepromCache_io_out_addr + io_gameConfig_eepromOffset[24:0]);
  assign _sdramArbiter_io_in_3_addr =
    25'(_soundRomCache_0_io_out_addr + io_gameConfig_sound_0_romOffset[24:0]);
  assign _sdramArbiter_io_in_4_addr =
    25'(_soundRomCache_1_io_out_addr + io_gameConfig_sound_1_romOffset[24:0]);
  assign _sdramArbiter_io_in_5_addr =
    25'(_layerRomCache_0_io_out_addr + io_gameConfig_layer_0_romOffset[24:0]);
  assign _sdramArbiter_io_in_6_addr =
    25'(_layerRomCache_1_io_out_addr + io_gameConfig_layer_1_romOffset[24:0]);
  assign _sdramArbiter_io_in_7_addr =
    25'(_layerRomCache_2_io_out_addr + io_gameConfig_layer_2_romOffset[24:0]);
  BurstMemArbiter_1 sdramArbiter (
    .clock             (clock),
    .reset             (reset),
    .io_in_0_wr        (_sdramDownloadBuffer_io_out_wr),
    .io_in_0_addr      (_sdramDownloadBuffer_io_out_addr),
    .io_in_0_din       (_sdramDownloadBuffer_io_out_din),
    .io_in_0_wait_n    (_sdramDownloadBuffer_io_out_wait_n),
    .io_in_0_burstDone (_sdramDownloadBuffer_io_out_burstDone),
    .io_in_1_rd        (_progRomCache_io_out_rd),
    .io_in_1_addr      (_progRomCache_io_out_addr),
    .io_in_1_dout      (_progRomCache_io_out_dout),
    .io_in_1_wait_n    (_progRomCache_io_out_wait_n),
    .io_in_1_valid     (_progRomCache_io_out_valid),
    .io_in_2_rd        (_eepromCache_io_out_rd),
    .io_in_2_wr        (_eepromCache_io_out_wr),
    .io_in_2_addr      (_sdramArbiter_io_in_2_addr),
    .io_in_2_din       (_eepromCache_io_out_din),
    .io_in_2_dout      (_eepromCache_io_out_dout),
    .io_in_2_wait_n    (_eepromCache_io_out_wait_n),
    .io_in_2_valid     (_eepromCache_io_out_valid),
    .io_in_3_rd        (_soundRomCache_0_io_out_rd),
    .io_in_3_addr      (_sdramArbiter_io_in_3_addr),
    .io_in_3_dout      (_soundRomCache_0_io_out_dout),
    .io_in_3_wait_n    (_soundRomCache_0_io_out_wait_n),
    .io_in_3_valid     (_soundRomCache_0_io_out_valid),
    .io_in_4_rd        (_soundRomCache_1_io_out_rd),
    .io_in_4_addr      (_sdramArbiter_io_in_4_addr),
    .io_in_4_dout      (_soundRomCache_1_io_out_dout),
    .io_in_4_wait_n    (_soundRomCache_1_io_out_wait_n),
    .io_in_4_valid     (_soundRomCache_1_io_out_valid),
    .io_in_5_rd        (_layerRomCache_0_io_out_rd),
    .io_in_5_addr      (_sdramArbiter_io_in_5_addr),
    .io_in_5_dout      (_layerRomCache_0_io_out_dout),
    .io_in_5_wait_n    (_layerRomCache_0_io_out_wait_n),
    .io_in_5_valid     (_layerRomCache_0_io_out_valid),
    .io_in_6_rd        (_layerRomCache_1_io_out_rd),
    .io_in_6_addr      (_sdramArbiter_io_in_6_addr),
    .io_in_6_dout      (_layerRomCache_1_io_out_dout),
    .io_in_6_wait_n    (_layerRomCache_1_io_out_wait_n),
    .io_in_6_valid     (_layerRomCache_1_io_out_valid),
    .io_in_7_rd        (_layerRomCache_2_io_out_rd),
    .io_in_7_addr      (_sdramArbiter_io_in_7_addr),
    .io_in_7_dout      (_layerRomCache_2_io_out_dout),
    .io_in_7_wait_n    (_layerRomCache_2_io_out_wait_n),
    .io_in_7_valid     (_layerRomCache_2_io_out_valid),
    .io_out_rd         (io_sdram_rd),
    .io_out_wr         (io_sdram_wr),
    .io_out_addr       (io_sdram_addr),
    .io_out_din        (io_sdram_din),
    .io_out_dout       (io_sdram_dout),
    .io_out_wait_n     (io_sdram_wait_n),
    .io_out_valid      (io_sdram_valid),
    .io_out_burstDone  (io_sdram_burstDone)
  );
  assign _nvramArbiter_io_in_0_addr = io_prog_nvram_addr[6:0];
  AsyncMemArbiter nvramArbiter (
    .clock          (clock),
    .reset          (reset),
    .io_in_0_rd     (io_prog_nvram_rd),
    .io_in_0_wr     (io_prog_nvram_wr),
    .io_in_0_addr   (_nvramArbiter_io_in_0_addr),
    .io_in_0_din    (io_prog_nvram_din),
    .io_in_0_dout   (io_prog_nvram_dout),
    .io_in_0_wait_n (io_prog_nvram_wait_n),
    .io_in_0_valid  (io_prog_nvram_valid),
    .io_in_1_rd     (io_eeprom_rd),
    .io_in_1_wr     (io_eeprom_wr),
    .io_in_1_addr   (io_eeprom_addr),
    .io_in_1_din    (io_eeprom_din),
    .io_in_1_dout   (io_eeprom_dout),
    .io_in_1_wait_n (io_eeprom_wait_n),
    .io_in_1_valid  (io_eeprom_valid),
    .io_out_rd      (_eepromCache_io_in_rd),
    .io_out_wr      (_eepromCache_io_in_wr),
    .io_out_addr    (_eepromCache_io_in_addr),
    .io_out_din     (_eepromCache_io_in_din),
    .io_out_dout    (_eepromCache_io_in_dout),
    .io_out_wait_n  (_eepromCache_io_in_wait_n),
    .io_out_valid   (_eepromCache_io_in_valid)
  );
  assign io_prog_rom_wait_n = _sdramDownloadBuffer_io_in_wait_n;
  assign io_ready = io_ready_enableReg;
endmodule

