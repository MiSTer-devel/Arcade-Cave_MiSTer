module TrueDualPortRam_11(
  input         clock,
  input         io_clockB,
  input         io_portA_wr,
  input  [6:0]  io_portA_addr,
  input  [63:0] io_portA_din,
  input  [8:0]  io_portB_addr,
  output [15:0] io_portB_dout
);

  wire       _ram_rd_a = 1'h0;
  wire [7:0] _ram_mask_a = 8'hFF;
  wire       _ram_rd_b = 1'h1;
  true_dual_port_ram #(
    .ADDR_WIDTH_A(7),
    .ADDR_WIDTH_B(9),
    .DATA_WIDTH_A(64),
    .DATA_WIDTH_B(16),
    .DEPTH_A(128),
    .DEPTH_B(512),
    .MASK_ENABLE("FALSE")
  ) ram (
    .clk_a  (clock),
    .rd_a   (_ram_rd_a),
    .wr_a   (io_portA_wr),
    .addr_a (io_portA_addr),
    .mask_a (_ram_mask_a),
    .din_a  (io_portA_din),
    .dout_a (/* unused */),
    .clk_b  (io_clockB),
    .rd_b   (_ram_rd_b),
    .addr_b (io_portB_addr),
    .dout_b (io_portB_dout)
  );
endmodule

